
module SME ( clk, reset, chardata, isstring, ispattern, valid, match, 
        match_index );
  input [7:0] chardata;
  output [4:0] match_index;
  input clk, reset, isstring, ispattern;
  output valid, match;
  wire   n4002, n4003, n4004, special, N166, N167, N168, N169, N170, N173,
         N174, N175, N176, N186, N187, N245, N246, N247, N842, N850, N851,
         N856, N857, N858, N1243, N1244, N1245, N1246, n374, n375, n449, n451,
         n452, n453, n589, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1709, n1711, n1713, n1715, n1717, n1719, n1720,
         n1721, n1722, n1723, N241, N240, N235, N234, N233,
         \add_802_S2/carry[5] , \add_802_S2/carry[4] , \add_802_S2/carry[3] ,
         \add_802_S2/carry[2] , \add_653_S2/carry[3] , \add_653_S2/carry[2] ,
         \add_653_S2/carry[1] , \r720/carry[4] , \r720/carry[3] ,
         \r720/carry[2] , \sub_1_root_sub_52_S2_2/carry[3] ,
         \sub_1_root_sub_52_S2_2/carry[2] , \sub_1_root_sub_52_S2_2/carry[1] ,
         \add_0_root_add_51/carry[5] , \add_0_root_add_51/carry[4] ,
         \add_0_root_add_51/carry[3] , \add_0_root_add_51/carry[2] , n3297,
         n6479, \r685/carry[2] , \r685/carry[3] , \r685/carry[4] ,
         \sub_1_root_add_0_root_add_92_2/n3 ,
         \sub_1_root_add_0_root_add_92_2/n1 ,
         \sub_1_root_add_0_root_add_92_2/carry[1] ,
         \sub_1_root_add_0_root_add_92_2/carry[2] ,
         \sub_1_root_add_0_root_add_92_2/carry[3] ,
         \sub_1_root_add_0_root_add_92_2/carry[4] ,
         \add_0_root_add_0_root_add_92_2/n1 ,
         \add_0_root_add_0_root_add_92_2/carry[2] ,
         \add_0_root_add_0_root_add_92_2/carry[3] ,
         \add_0_root_add_0_root_add_92_2/carry[4] , n6478, n4426, n4427, n4428,
         n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438,
         n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448,
         n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458,
         n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468,
         n4469, n4470, n4471, n4473, n4474, n4475, n4477, n4478, n4490, n4492,
         n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
         n4515, n4516, n4518, n4527, n4537, n4538, n4542, n4544, n4545, n4546,
         n4547, n4548, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4561,
         n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571,
         n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581,
         n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591,
         n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601,
         n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611,
         n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621,
         n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631,
         n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641,
         n4642, n4643, n4648, n4649, n4652, n4653, n4654, n4655, n4656, n4657,
         n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668,
         n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678,
         n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688,
         n4689, n4690, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699,
         n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709,
         n4710, n4711, n4712, n4713, n4715, n4716, n4717, n4718, n4719, n4720,
         n4721, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731,
         n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741,
         n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751,
         n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4832, n4833,
         n4834, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844,
         n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854,
         n4855, n4856, n4857, n4858, n4859, n4860, n4863, n4867, n4868, n4869,
         n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4911,
         n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921,
         n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931,
         n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941,
         n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951,
         n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961,
         n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971,
         n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981,
         n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991,
         n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001,
         n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011,
         n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021,
         n5022, n5023, n5024, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5330, n5331, n5332, n5333,
         n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343,
         n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353,
         n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363,
         n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373,
         n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383,
         n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393,
         n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403,
         n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413,
         n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423,
         n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433,
         n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443,
         n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453,
         n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463,
         n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473,
         n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483,
         n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493,
         n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503,
         n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513,
         n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523,
         n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533,
         n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543,
         n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553,
         n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563,
         n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573,
         n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583,
         n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593,
         n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603,
         n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613,
         n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623,
         n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633,
         n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643,
         n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653,
         n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663,
         n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673,
         n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683,
         n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693,
         n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5704,
         n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714,
         n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724,
         n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734,
         n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744,
         n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754,
         n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764,
         n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774,
         n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784,
         n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794,
         n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804,
         n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814,
         n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824,
         n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834,
         n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844,
         n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854,
         n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864,
         n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874,
         n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884,
         n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894,
         n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904,
         n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914,
         n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924,
         n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934,
         n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944,
         n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954,
         n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5968, n5969,
         n5970, n5971, n5972, n5973, n5974, n5975, n5977, n5978, n5979, n5980,
         n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990,
         n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000,
         n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010,
         n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020,
         n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030,
         n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040,
         n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050,
         n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060,
         n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070,
         n6071, n6073, n6074, n6075, n6275, n6276, n6277, n6278, n6279, n6280,
         n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290,
         n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300,
         n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310,
         n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320,
         n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330,
         n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340,
         n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350,
         n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360,
         n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370,
         n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380,
         n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390,
         n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400,
         n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410,
         n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420,
         n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430,
         n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440,
         n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450,
         n6451, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6471, n6472, n6473,
         n6474, n6476, n6477;
  wire   [5:0] stringNum;
  wire   [3:0] patternCounter;
  wire   [63:0] pattern;
  wire   [2:0] special_locate;
  wire   [2:0] next_state;
  wire   [255:0] stringData;
  wire   [63:0] pattern_after;
  wire   [5:0] stringCounter;

  OAI31X2 U3220 ( .A0(n4997), .A1(n6348), .A2(n4834), .B0(n4989), .Y(n4999) );
  OAI31X2 U3322 ( .A0(n5034), .A1(n5035), .A2(n5036), .B0(n6308), .Y(n5026) );
  OAI31X2 U3326 ( .A0(n6290), .A1(n5034), .A2(n4544), .B0(n6308), .Y(n5019) );
  OAI221X2 U3343 ( .A0(n4857), .A1(n5042), .B0(n5043), .B1(n5016), .C0(n5044), 
        .Y(next_state[2]) );
  OAI221X2 U3345 ( .A0(special), .A1(n5042), .B0(n4470), .B1(n5016), .C0(n5046), .Y(next_state[1]) );
  OAI211X2 U3365 ( .A0(n5063), .A1(n4468), .B0(n5064), .C0(n5016), .Y(
        next_state[0]) );
  OAI221X2 U3896 ( .A0(n5017), .A1(n4686), .B0(n6457), .B1(n5696), .C0(n5697), 
        .Y(n5355) );
  OAI221X2 U3906 ( .A0(n5017), .A1(n4689), .B0(n6457), .B1(n5709), .C0(n5710), 
        .Y(n5364) );
  OAI221X2 U3911 ( .A0(n5017), .A1(n4687), .B0(n6457), .B1(n5713), .C0(n5714), 
        .Y(n5360) );
  DFFRX1 \matc_indexTemp_reg[3]  ( .D(n1374), .CK(clk), .RN(n6427), .QN(n5958)
         );
  DFFRX1 \matc_indexTemp_reg[1]  ( .D(n1378), .CK(clk), .RN(n6427), .QN(n5961)
         );
  DFFRX1 \matc_indexTemp_reg[2]  ( .D(n1376), .CK(clk), .RN(n6426), .QN(n5959)
         );
  DFFRX1 \matc_indexTemp_reg[4]  ( .D(n1721), .CK(clk), .RN(n6427), .QN(n5960)
         );
  DFFRX1 \matc_indexTemp_reg[0]  ( .D(n1380), .CK(clk), .RN(n6427), .QN(n5962)
         );
  DFFRX1 \current_state_reg[0]  ( .D(n6276), .CK(clk), .RN(n6421), .QN(n375)
         );
  DFFRX1 \pattern_after_reg[48]  ( .D(n1367), .CK(clk), .RN(n6431), .QN(n6052)
         );
  DFFRX1 \pattern_after_reg[50]  ( .D(n1353), .CK(clk), .RN(n6432), .Q(
        pattern_after[50]), .QN(n6069) );
  DFFRX1 \pattern_after_reg[42]  ( .D(n1354), .CK(clk), .RN(n6432), .Q(
        pattern_after[42]), .QN(n6064) );
  DFFRX1 \pattern_after_reg[53]  ( .D(n1337), .CK(clk), .RN(n6432), .Q(
        pattern_after[53]), .QN(n6068) );
  DFFRX1 \pattern_after_reg[45]  ( .D(n1332), .CK(clk), .RN(n6432), .Q(
        pattern_after[45]), .QN(n6062) );
  DFFRX1 \pattern_after_reg[49]  ( .D(n1365), .CK(clk), .RN(n6431), .Q(
        pattern_after[49]), .QN(n6060) );
  DFFRX1 \pattern_after_reg[41]  ( .D(n1360), .CK(clk), .RN(n6431), .Q(
        pattern_after[41]), .QN(n6001) );
  DFFRX1 \pattern_after_reg[33]  ( .D(n1361), .CK(clk), .RN(n6430), .Q(
        pattern_after[33]), .QN(n5998) );
  DFFRX1 \pattern_after_reg[51]  ( .D(n1351), .CK(clk), .RN(n6431), .Q(
        pattern_after[51]), .QN(n6005) );
  DFFRX1 \pattern_after_reg[43]  ( .D(n1346), .CK(clk), .RN(n6431), .Q(
        pattern_after[43]), .QN(n6053) );
  DFFRX1 \pattern_after_reg[35]  ( .D(n1347), .CK(clk), .RN(n6424), .Q(
        pattern_after[35]), .QN(n6043) );
  DFFRX1 \pattern_after_reg[55]  ( .D(n1323), .CK(clk), .RN(n6431), .Q(
        pattern_after[55]), .QN(n6066) );
  DFFRX1 \pattern_after_reg[52]  ( .D(n1344), .CK(clk), .RN(n6431), .Q(
        pattern_after[52]), .QN(n6067) );
  DFFRX1 \pattern_after_reg[54]  ( .D(n1330), .CK(clk), .RN(n6431), .Q(
        pattern_after[54]) );
  DFFRX1 \pattern_after_reg[34]  ( .D(n1355), .CK(clk), .RN(n6431), .Q(
        pattern_after[34]), .QN(n6058) );
  DFFRX1 \pattern_after_reg[26]  ( .D(n1356), .CK(clk), .RN(n6431), .Q(
        pattern_after[26]), .QN(n6050) );
  DFFRX1 \pattern_after_reg[29]  ( .D(n1334), .CK(clk), .RN(n6431), .Q(
        pattern_after[29]), .QN(n6049) );
  DFFRX1 \pattern_after_reg[37]  ( .D(n1333), .CK(clk), .RN(n6416), .Q(
        pattern_after[37]), .QN(n6057) );
  DFFRX1 \pattern_after_reg[32]  ( .D(n1369), .CK(clk), .RN(n6430), .Q(n5974), 
        .QN(n5995) );
  DFFRX1 \pattern_after_reg[24]  ( .D(n1370), .CK(clk), .RN(n6430), .Q(n5975), 
        .QN(n5993) );
  DFFRX1 \pattern_after_reg[40]  ( .D(n1368), .CK(clk), .RN(n6431), .Q(n5973), 
        .QN(n5999) );
  DFFRX1 \pattern_after_reg[8]  ( .D(n1372), .CK(clk), .RN(n6417), .Q(
        pattern_after[8]), .QN(n5981) );
  DFFRX1 \pattern_after_reg[14]  ( .D(n1329), .CK(clk), .RN(n6417), .Q(
        pattern_after[14]), .QN(n5979) );
  DFFRX1 \pattern_after_reg[25]  ( .D(n1362), .CK(clk), .RN(n6430), .Q(
        pattern_after[25]), .QN(n5994) );
  DFFRX1 \pattern_after_reg[17]  ( .D(n1363), .CK(clk), .RN(n6418), .Q(
        pattern_after[17]), .QN(n5992) );
  DFFRX1 \pattern_after_reg[27]  ( .D(n1348), .CK(clk), .RN(n6430), .Q(
        pattern_after[27]), .QN(n6036) );
  DFFRX1 \pattern_after_reg[19]  ( .D(n1349), .CK(clk), .RN(n6418), .Q(
        pattern_after[19]), .QN(n6035) );
  DFFRX1 \pattern_after_reg[12]  ( .D(n1343), .CK(clk), .RN(n6417), .Q(
        pattern_after[12]), .QN(n5996) );
  DFFRX1 \pattern_after_reg[15]  ( .D(n1322), .CK(clk), .RN(n6418), .Q(
        pattern_after[15]), .QN(n6037) );
  DFFRX1 \pattern_after_reg[47]  ( .D(n1318), .CK(clk), .RN(n6430), .Q(
        pattern_after[47]), .QN(n6054) );
  DFFRX1 \pattern_after_reg[46]  ( .D(n1325), .CK(clk), .RN(n6430), .Q(
        pattern_after[46]), .QN(n6002) );
  DFFRX1 \pattern_after_reg[28]  ( .D(n1341), .CK(clk), .RN(n6430), .Q(
        pattern_after[28]), .QN(n6038) );
  DFFRX1 \pattern_after_reg[36]  ( .D(n1340), .CK(clk), .RN(n6420), .Q(
        pattern_after[36]), .QN(n6044) );
  DFFRX1 \pattern_after_reg[39]  ( .D(n1319), .CK(clk), .RN(n6416), .Q(
        pattern_after[39]), .QN(n6003) );
  DFFRX1 \pattern_after_reg[30]  ( .D(n1327), .CK(clk), .RN(n6430), .Q(
        pattern_after[30]), .QN(n6045) );
  DFFRX1 \pattern_after_reg[31]  ( .D(n1320), .CK(clk), .RN(n6430), .Q(
        pattern_after[31]), .QN(n6000) );
  DFFRX1 \pattern_after_reg[38]  ( .D(n1326), .CK(clk), .RN(n6416), .Q(
        pattern_after[38]), .QN(n6055) );
  DFFRX1 \pattern_after_reg[44]  ( .D(n1339), .CK(clk), .RN(n6430), .Q(
        pattern_after[44]), .QN(n6061) );
  EDFFX1 \stringNum_reg[5]  ( .D(stringCounter[5]), .E(n3297), .CK(clk), .Q(
        stringNum[5]) );
  DFFRX1 \pattern_after_reg[18]  ( .D(n1357), .CK(clk), .RN(n6418), .Q(
        pattern_after[18]), .QN(n6042) );
  DFFRX1 \pattern_after_reg[21]  ( .D(n1335), .CK(clk), .RN(n6418), .Q(
        pattern_after[21]), .QN(n6041) );
  DFFRX1 \pattern_after_reg[16]  ( .D(n1371), .CK(clk), .RN(n6428), .Q(n5972), 
        .QN(n5990) );
  DFFRX1 \pattern_after_reg[9]  ( .D(n1364), .CK(clk), .RN(n6427), .Q(n5968)
         );
  DFFRX1 \pattern_after_reg[13]  ( .D(n1336), .CK(clk), .RN(n6428), .Q(n5969)
         );
  DFFRX1 \pattern_after_reg[11]  ( .D(n1350), .CK(clk), .RN(n6428), .Q(n5970)
         );
  DFFRX1 \pattern_after_reg[10]  ( .D(n1358), .CK(clk), .RN(n6428), .Q(n5971)
         );
  DFFRX1 \special_locate_reg[0]  ( .D(n1451), .CK(clk), .RN(n6427), .Q(n5991), 
        .QN(n589) );
  DFFRX1 \pattern_after_reg[22]  ( .D(n1328), .CK(clk), .RN(n6418), .Q(
        pattern_after[22]), .QN(n6039) );
  DFFRX1 \pattern_after_reg[20]  ( .D(n1342), .CK(clk), .RN(n6418), .Q(
        pattern_after[20]), .QN(n5997) );
  EDFFX1 \stringNum_reg[2]  ( .D(stringCounter[2]), .E(n3297), .CK(clk), .Q(
        stringNum[2]) );
  EDFFX1 \stringNum_reg[1]  ( .D(stringCounter[1]), .E(n3297), .CK(clk), .Q(
        stringNum[1]) );
  DFFRX1 \pattern_after_reg[23]  ( .D(n1321), .CK(clk), .RN(n6418), .Q(
        pattern_after[23]), .QN(n6040) );
  DFFRX1 \pattern_reg[58]  ( .D(n1387), .CK(clk), .RN(n6429), .Q(pattern[58]), 
        .QN(n6070) );
  DFFRX1 \pattern_reg[50]  ( .D(n1395), .CK(clk), .RN(n6429), .Q(pattern[50]), 
        .QN(n6065) );
  DFFRX1 \pattern_reg[42]  ( .D(n1403), .CK(clk), .RN(n6429), .Q(pattern[42]), 
        .QN(n6059) );
  DFFRX1 \pattern_reg[34]  ( .D(n1411), .CK(clk), .RN(n6429), .Q(pattern[34]), 
        .QN(n6051) );
  DFFRX1 \pattern_after_reg[3]  ( .D(n1352), .CK(clk), .RN(n6418), .Q(
        pattern_after[3]), .QN(n6034) );
  DFFRX1 \pattern_after_reg[2]  ( .D(n1359), .CK(clk), .RN(n6418), .Q(
        pattern_after[2]), .QN(n6032) );
  DFFRX1 \pattern_reg[61]  ( .D(n1384), .CK(clk), .RN(n6429), .Q(pattern[61]), 
        .QN(n6063) );
  DFFRX1 \pattern_reg[53]  ( .D(n1392), .CK(clk), .RN(n6429), .Q(pattern[53]), 
        .QN(n6056) );
  DFFRX1 \pattern_reg[45]  ( .D(n1400), .CK(clk), .RN(n6429), .Q(pattern[45]), 
        .QN(n6048) );
  DFFRX1 \pattern_reg[37]  ( .D(n1408), .CK(clk), .RN(n6428), .Q(pattern[37]), 
        .QN(n6047) );
  DFFRX1 \pattern_after_reg[1]  ( .D(n1366), .CK(clk), .RN(n6418), .Q(
        pattern_after[1]), .QN(n6033) );
  DFFRX1 \pattern_reg[56]  ( .D(n1389), .CK(clk), .RN(n6428), .Q(pattern[56]), 
        .QN(n6017) );
  DFFRX1 \pattern_reg[48]  ( .D(n1397), .CK(clk), .RN(n6428), .Q(pattern[48]), 
        .QN(n6020) );
  DFFRX1 \pattern_reg[40]  ( .D(n1405), .CK(clk), .RN(n6428), .Q(pattern[40]), 
        .QN(n6019) );
  DFFRX1 \pattern_reg[32]  ( .D(n1413), .CK(clk), .RN(n6428), .Q(pattern[32]), 
        .QN(n6018) );
  DFFRX1 \pattern_after_reg[6]  ( .D(n1331), .CK(clk), .RN(n6419), .Q(
        pattern_after[6]), .QN(n5985) );
  DFFRX1 \pattern_after_reg[5]  ( .D(n1338), .CK(clk), .RN(n6419), .Q(
        pattern_after[5]), .QN(n6014) );
  DFFRX1 \pattern_after_reg[4]  ( .D(n1345), .CK(clk), .RN(n6419), .Q(
        pattern_after[4]), .QN(n6013) );
  DFFRX1 \pattern_reg[57]  ( .D(n1388), .CK(clk), .RN(n6430), .Q(pattern[57]), 
        .QN(n6026) );
  DFFRX1 \pattern_reg[49]  ( .D(n1396), .CK(clk), .RN(n6429), .Q(pattern[49]), 
        .QN(n6025) );
  DFFRX1 \pattern_reg[41]  ( .D(n1404), .CK(clk), .RN(n6429), .Q(pattern[41]), 
        .QN(n6024) );
  DFFRX1 \pattern_reg[33]  ( .D(n1412), .CK(clk), .RN(n6428), .Q(pattern[33]), 
        .QN(n6023) );
  DFFRX1 \pattern_reg[59]  ( .D(n1386), .CK(clk), .RN(n6429), .Q(pattern[59]), 
        .QN(n5989) );
  DFFRX1 \pattern_reg[51]  ( .D(n1394), .CK(clk), .RN(n6429), .Q(pattern[51]), 
        .QN(n5987) );
  DFFRX1 \pattern_reg[43]  ( .D(n1402), .CK(clk), .RN(n6429), .Q(pattern[43]), 
        .QN(n5988) );
  DFFRX1 \pattern_reg[35]  ( .D(n1410), .CK(clk), .RN(n6428), .Q(pattern[35]), 
        .QN(n5986) );
  DFFRX1 \pattern_reg[63]  ( .D(n1382), .CK(clk), .RN(n6423), .Q(pattern[63])
         );
  DFFRX1 \pattern_reg[47]  ( .D(n1398), .CK(clk), .RN(n6422), .Q(pattern[47])
         );
  DFFRX1 \pattern_reg[39]  ( .D(n1406), .CK(clk), .RN(n6422), .Q(pattern[39])
         );
  DFFRX1 \pattern_reg[55]  ( .D(n1390), .CK(clk), .RN(n6422), .Q(pattern[55])
         );
  DFFRX1 \pattern_reg[62]  ( .D(n1383), .CK(clk), .RN(n6422), .Q(pattern[62])
         );
  DFFRX1 \pattern_reg[46]  ( .D(n1399), .CK(clk), .RN(n6422), .Q(pattern[46])
         );
  DFFRX1 \pattern_reg[38]  ( .D(n1407), .CK(clk), .RN(n6422), .Q(pattern[38])
         );
  DFFRX1 \pattern_reg[54]  ( .D(n1391), .CK(clk), .RN(n6422), .Q(pattern[54])
         );
  DFFRX1 \pattern_reg[60]  ( .D(n1385), .CK(clk), .RN(n6422), .Q(pattern[60])
         );
  DFFRX1 \pattern_reg[44]  ( .D(n1401), .CK(clk), .RN(n6422), .Q(pattern[44])
         );
  DFFRX1 \pattern_reg[36]  ( .D(n1409), .CK(clk), .RN(n6422), .Q(pattern[36])
         );
  DFFRX1 \pattern_reg[52]  ( .D(n1393), .CK(clk), .RN(n6422), .Q(pattern[52])
         );
  DFFRX1 \pattern_after_reg[7]  ( .D(n1324), .CK(clk), .RN(n6419), .Q(
        pattern_after[7]) );
  DFFRX1 \pattern_after_reg[0]  ( .D(n1373), .CK(clk), .RN(n6418), .Q(
        pattern_after[0]) );
  DFFRX1 \pattern_reg[10]  ( .D(n1435), .CK(clk), .RN(n6427), .QN(n5978) );
  DFFRX1 \pattern_reg[11]  ( .D(n1434), .CK(clk), .RN(n6427), .QN(n5984) );
  DFFRX1 \pattern_reg[13]  ( .D(n1432), .CK(clk), .RN(n6427), .QN(n5980) );
  DFFRX1 \pattern_reg[9]  ( .D(n1436), .CK(clk), .RN(n6427), .QN(n6011) );
  DFFRX1 \stringData_reg[129]  ( .D(n1578), .CK(clk), .RN(n6414), .QN(n6012)
         );
  DFFRX1 \stringData_reg[31]  ( .D(n1676), .CK(clk), .RN(n6434), .Q(
        stringData[31]) );
  DFFRX1 \stringData_reg[30]  ( .D(n1677), .CK(clk), .RN(n6434), .Q(
        stringData[30]) );
  DFFRX1 \stringData_reg[29]  ( .D(n1678), .CK(clk), .RN(n6434), .Q(
        stringData[29]) );
  DFFRX1 \stringData_reg[28]  ( .D(n1679), .CK(clk), .RN(n6434), .Q(
        stringData[28]) );
  DFFRX1 \stringData_reg[27]  ( .D(n1680), .CK(clk), .RN(n6433), .Q(
        stringData[27]) );
  DFFRX1 \stringData_reg[26]  ( .D(n1681), .CK(clk), .RN(n6433), .Q(
        stringData[26]) );
  DFFRX1 \stringData_reg[25]  ( .D(n1682), .CK(clk), .RN(n6433), .Q(
        stringData[25]) );
  DFFRX1 \stringData_reg[24]  ( .D(n1683), .CK(clk), .RN(n6433), .Q(
        stringData[24]) );
  DFFRX1 \stringData_reg[23]  ( .D(n1684), .CK(clk), .RN(n6433), .Q(
        stringData[23]) );
  DFFRX1 \stringData_reg[22]  ( .D(n1685), .CK(clk), .RN(n6433), .Q(
        stringData[22]) );
  DFFRX1 \stringData_reg[21]  ( .D(n1686), .CK(clk), .RN(n6433), .Q(
        stringData[21]) );
  DFFRX1 \stringData_reg[20]  ( .D(n1687), .CK(clk), .RN(n6433), .Q(
        stringData[20]) );
  DFFRX1 \stringData_reg[19]  ( .D(n1688), .CK(clk), .RN(n6433), .Q(
        stringData[19]) );
  DFFRX1 \stringData_reg[18]  ( .D(n1689), .CK(clk), .RN(n6433), .Q(
        stringData[18]) );
  DFFRX1 \stringData_reg[17]  ( .D(n1690), .CK(clk), .RN(n6433), .Q(
        stringData[17]) );
  DFFRX1 \stringData_reg[16]  ( .D(n1691), .CK(clk), .RN(n6433), .Q(
        stringData[16]) );
  DFFRX1 \stringData_reg[39]  ( .D(n1668), .CK(clk), .RN(n6438), .Q(
        stringData[39]) );
  DFFRX1 \stringData_reg[38]  ( .D(n1669), .CK(clk), .RN(n6438), .Q(
        stringData[38]) );
  DFFRX1 \stringData_reg[37]  ( .D(n1670), .CK(clk), .RN(n6438), .Q(
        stringData[37]) );
  DFFRX1 \stringData_reg[36]  ( .D(n1671), .CK(clk), .RN(n6438), .Q(
        stringData[36]) );
  DFFRX1 \stringData_reg[35]  ( .D(n1672), .CK(clk), .RN(n6438), .Q(
        stringData[35]) );
  DFFRX1 \stringData_reg[34]  ( .D(n1673), .CK(clk), .RN(n6437), .Q(
        stringData[34]) );
  DFFRX1 \stringData_reg[33]  ( .D(n1674), .CK(clk), .RN(n6437), .Q(
        stringData[33]) );
  DFFRX1 \stringData_reg[32]  ( .D(n1675), .CK(clk), .RN(n6437), .Q(
        stringData[32]) );
  DFFRX1 \stringData_reg[119]  ( .D(n1588), .CK(clk), .RN(n6435), .Q(
        stringData[119]), .QN(n6007) );
  DFFRX1 \pattern_reg[3]  ( .D(n1442), .CK(clk), .RN(n6417), .Q(pattern[3]), 
        .QN(n6016) );
  DFFRX1 \pattern_reg[2]  ( .D(n1443), .CK(clk), .RN(n6416), .Q(pattern[2]), 
        .QN(n6031) );
  DFFRX1 \stringData_reg[255]  ( .D(n1452), .CK(clk), .RN(n6424), .Q(
        stringData[255]) );
  DFFRX1 \stringData_reg[253]  ( .D(n1454), .CK(clk), .RN(n6424), .Q(
        stringData[253]) );
  DFFRX1 \stringData_reg[250]  ( .D(n1457), .CK(clk), .RN(n6424), .Q(
        stringData[250]) );
  DFFRX1 \stringData_reg[248]  ( .D(n1459), .CK(clk), .RN(n6424), .Q(
        stringData[248]) );
  DFFRX1 \stringData_reg[15]  ( .D(n1692), .CK(clk), .RN(n6437), .Q(
        stringData[15]) );
  DFFRX1 \stringData_reg[14]  ( .D(n1693), .CK(clk), .RN(n6437), .Q(
        stringData[14]) );
  DFFRX1 \stringData_reg[13]  ( .D(n1694), .CK(clk), .RN(n6437), .Q(
        stringData[13]) );
  DFFRX1 \stringData_reg[12]  ( .D(n1695), .CK(clk), .RN(n6437), .Q(
        stringData[12]) );
  DFFRX1 \stringData_reg[11]  ( .D(n1696), .CK(clk), .RN(n6437), .Q(
        stringData[11]) );
  DFFRX1 \stringData_reg[10]  ( .D(n1697), .CK(clk), .RN(n6437), .Q(
        stringData[10]) );
  DFFRX1 \stringData_reg[9]  ( .D(n1698), .CK(clk), .RN(n6437), .Q(
        stringData[9]) );
  DFFRX1 \stringData_reg[8]  ( .D(n1699), .CK(clk), .RN(n6437), .Q(
        stringData[8]) );
  DFFRX1 \stringData_reg[127]  ( .D(n1580), .CK(clk), .RN(n6436), .Q(
        stringData[127]) );
  DFFRX1 \stringData_reg[125]  ( .D(n1582), .CK(clk), .RN(n6436), .Q(
        stringData[125]) );
  DFFRX1 \stringData_reg[122]  ( .D(n1585), .CK(clk), .RN(n6435), .Q(
        stringData[122]) );
  DFFRX1 \stringData_reg[120]  ( .D(n1587), .CK(clk), .RN(n6435), .Q(
        stringData[120]) );
  DFFRX1 \pattern_reg[1]  ( .D(n1444), .CK(clk), .RN(n6416), .Q(pattern[1]), 
        .QN(n6015) );
  DFFRX1 \stringData_reg[105]  ( .D(n1602), .CK(clk), .RN(n6426), .Q(
        stringData[105]), .QN(n6046) );
  DFFRX1 \pattern_reg[6]  ( .D(n1439), .CK(clk), .RN(n6417), .Q(pattern[6]), 
        .QN(n5983) );
  DFFRX1 \pattern_reg[5]  ( .D(n1440), .CK(clk), .RN(n6417), .Q(pattern[5]), 
        .QN(n6008) );
  DFFRX1 \pattern_reg[4]  ( .D(n1441), .CK(clk), .RN(n6417), .Q(pattern[4]), 
        .QN(n6010) );
  DFFRX1 \pattern_reg[8]  ( .D(n1437), .CK(clk), .RN(n6417), .Q(pattern[8]), 
        .QN(n6027) );
  DFFRX1 \pattern_reg[15]  ( .D(n1430), .CK(clk), .RN(n6417), .Q(pattern[15]), 
        .QN(n6029) );
  DFFRX1 \pattern_reg[14]  ( .D(n1431), .CK(clk), .RN(n6417), .Q(pattern[14]), 
        .QN(n6028) );
  DFFRX1 \pattern_reg[12]  ( .D(n1433), .CK(clk), .RN(n6417), .Q(pattern[12]), 
        .QN(n6030) );
  DFFRX1 \stringData_reg[103]  ( .D(n1604), .CK(clk), .RN(n6426), .Q(
        stringData[103]) );
  DFFRX1 \stringData_reg[102]  ( .D(n1605), .CK(clk), .RN(n6426), .Q(
        stringData[102]) );
  DFFRX1 \stringData_reg[101]  ( .D(n1606), .CK(clk), .RN(n6426), .Q(
        stringData[101]) );
  DFFRX1 \stringData_reg[100]  ( .D(n1607), .CK(clk), .RN(n6425), .Q(
        stringData[100]) );
  DFFRX1 \stringData_reg[99]  ( .D(n1608), .CK(clk), .RN(n6425), .Q(
        stringData[99]) );
  DFFRX1 \stringData_reg[98]  ( .D(n1609), .CK(clk), .RN(n6425), .Q(
        stringData[98]) );
  DFFRX1 \stringData_reg[97]  ( .D(n1610), .CK(clk), .RN(n6425), .Q(
        stringData[97]) );
  DFFRX1 \stringData_reg[96]  ( .D(n1611), .CK(clk), .RN(n6425), .Q(
        stringData[96]) );
  DFFRX1 \stringData_reg[245]  ( .D(n1462), .CK(clk), .RN(n6423), .Q(
        stringData[245]) );
  DFFRX1 \stringData_reg[242]  ( .D(n1465), .CK(clk), .RN(n6423), .Q(
        stringData[242]) );
  DFFRX1 \stringData_reg[240]  ( .D(n1467), .CK(clk), .RN(n6423), .Q(
        stringData[240]) );
  DFFRX1 \stringData_reg[117]  ( .D(n1590), .CK(clk), .RN(n6435), .Q(
        stringData[117]) );
  DFFRX1 \stringData_reg[114]  ( .D(n1593), .CK(clk), .RN(n6435), .Q(
        stringData[114]) );
  DFFRX1 \stringData_reg[112]  ( .D(n1595), .CK(clk), .RN(n6435), .Q(
        stringData[112]) );
  DFFRX1 \stringData_reg[247]  ( .D(n1460), .CK(clk), .RN(n6423), .Q(
        stringData[247]) );
  DFFRX1 \stringData_reg[143]  ( .D(n1564), .CK(clk), .RN(n6415), .Q(
        stringData[143]) );
  DFFRX1 \stringData_reg[142]  ( .D(n1565), .CK(clk), .RN(n6415), .Q(
        stringData[142]) );
  DFFRX1 \stringData_reg[141]  ( .D(n1566), .CK(clk), .RN(n6415), .Q(
        stringData[141]) );
  DFFRX1 \stringData_reg[140]  ( .D(n1567), .CK(clk), .RN(n6415), .Q(
        stringData[140]) );
  DFFRX1 \stringData_reg[139]  ( .D(n1568), .CK(clk), .RN(n6415), .Q(
        stringData[139]) );
  DFFRX1 \stringData_reg[138]  ( .D(n1569), .CK(clk), .RN(n6415), .Q(
        stringData[138]) );
  DFFRX1 \stringData_reg[137]  ( .D(n1570), .CK(clk), .RN(n6415), .Q(
        stringData[137]) );
  DFFRX1 \stringData_reg[136]  ( .D(n1571), .CK(clk), .RN(n6414), .Q(
        stringData[136]) );
  DFFRX1 \stringData_reg[57]  ( .D(n1650), .CK(clk), .RN(n6075), .QN(n5982) );
  DFFRX1 \stringData_reg[49]  ( .D(n1658), .CK(clk), .RN(n6434), .QN(n6009) );
  DFFRX1 \stringData_reg[254]  ( .D(n1453), .CK(clk), .RN(n6424), .Q(
        stringData[254]) );
  DFFRX1 \stringData_reg[252]  ( .D(n1455), .CK(clk), .RN(n6424), .Q(
        stringData[252]) );
  DFFRX1 \stringData_reg[251]  ( .D(n1456), .CK(clk), .RN(n6424), .Q(
        stringData[251]) );
  DFFRX1 \stringData_reg[249]  ( .D(n1458), .CK(clk), .RN(n6424), .Q(
        stringData[249]) );
  DFFRX1 \stringData_reg[126]  ( .D(n1581), .CK(clk), .RN(n6436), .Q(
        stringData[126]) );
  DFFRX1 \stringData_reg[124]  ( .D(n1583), .CK(clk), .RN(n6436), .Q(
        stringData[124]) );
  DFFRX1 \stringData_reg[123]  ( .D(n1584), .CK(clk), .RN(n6436), .Q(
        stringData[123]) );
  DFFRX1 \stringData_reg[121]  ( .D(n1586), .CK(clk), .RN(n6435), .Q(
        stringData[121]) );
  DFFRX1 \match_index_reg[0]  ( .D(n1381), .CK(clk), .RN(n6420), .Q(n6479), 
        .QN(n6022) );
  DFFRX1 \stringData_reg[246]  ( .D(n1461), .CK(clk), .RN(n6423), .Q(
        stringData[246]) );
  DFFRX1 \stringData_reg[244]  ( .D(n1463), .CK(clk), .RN(n6423), .Q(
        stringData[244]) );
  DFFRX1 \stringData_reg[243]  ( .D(n1464), .CK(clk), .RN(n6423), .Q(
        stringData[243]) );
  DFFRX1 \stringData_reg[241]  ( .D(n1466), .CK(clk), .RN(n6423), .Q(
        stringData[241]) );
  DFFRX1 \stringData_reg[118]  ( .D(n1589), .CK(clk), .RN(n6435), .Q(
        stringData[118]) );
  DFFRX1 \stringData_reg[116]  ( .D(n1591), .CK(clk), .RN(n6435), .Q(
        stringData[116]) );
  DFFRX1 \stringData_reg[115]  ( .D(n1592), .CK(clk), .RN(n6435), .Q(
        stringData[115]) );
  DFFRX1 \stringData_reg[113]  ( .D(n1594), .CK(clk), .RN(n6435), .Q(
        stringData[113]) );
  ADDHXL U4688 ( .A(stringCounter[1]), .B(stringCounter[0]), .CO(
        \add_802_S2/carry[2] ), .S(N1243) );
  ADDHXL U4689 ( .A(stringCounter[3]), .B(\add_802_S2/carry[3] ), .CO(
        \add_802_S2/carry[4] ), .S(N1245) );
  ADDHXL U4690 ( .A(stringCounter[2]), .B(\add_802_S2/carry[2] ), .CO(
        \add_802_S2/carry[3] ), .S(N1244) );
  ADDHXL U4691 ( .A(stringCounter[4]), .B(\add_802_S2/carry[4] ), .CO(
        \add_802_S2/carry[5] ), .S(N1246) );
  ADDFXL U4683 ( .A(n4004), .B(special_locate[1]), .CI(\add_653_S2/carry[1] ), 
        .CO(\add_653_S2/carry[2] ), .S(N850) );
  ADDHXL U3863 ( .A(n4003), .B(\r720/carry[2] ), .CO(\r720/carry[3] ), .S(N857) );
  ADDHXL U3862 ( .A(n4004), .B(match_index[0]), .CO(\r720/carry[2] ), .S(N856)
         );
  ADDHXL U3864 ( .A(n4002), .B(\r720/carry[3] ), .CO(\r720/carry[4] ), .S(N858) );
  ADDFXL \add_0_root_add_0_root_add_92_2/U1_1  ( .A(n4859), .B(N233), .CI(
        \add_0_root_add_0_root_add_92_2/n1 ), .CO(
        \add_0_root_add_0_root_add_92_2/carry[2] ), .S(N245) );
  ADDFXL \add_0_root_add_0_root_add_92_2/U1_2  ( .A(N240), .B(N234), .CI(
        \add_0_root_add_0_root_add_92_2/carry[2] ), .CO(
        \add_0_root_add_0_root_add_92_2/carry[3] ), .S(N246) );
  ADDFXL \sub_1_root_add_0_root_add_92_2/U2_2  ( .A(stringNum[2]), .B(n4860), 
        .CI(\sub_1_root_add_0_root_add_92_2/carry[2] ), .CO(
        \sub_1_root_add_0_root_add_92_2/carry[3] ), .S(N234) );
  ADDFXL \sub_1_root_add_0_root_add_92_2/U2_1  ( .A(stringNum[1]), .B(n4834), 
        .CI(\sub_1_root_add_0_root_add_92_2/carry[1] ), .CO(
        \sub_1_root_add_0_root_add_92_2/carry[2] ), .S(N233) );
  ADDFXL \sub_1_root_add_0_root_add_92_2/U2_3  ( .A(stringNum[3]), .B(n6021), 
        .CI(\sub_1_root_add_0_root_add_92_2/carry[3] ), .CO(
        \sub_1_root_add_0_root_add_92_2/carry[4] ), .S(N235) );
  ADDFXL U4615 ( .A(stringNum[2]), .B(n4858), .CI(
        \sub_1_root_sub_52_S2_2/carry[2] ), .CO(
        \sub_1_root_sub_52_S2_2/carry[3] ), .S(N187) );
  ADDFXL U4617 ( .A(stringNum[1]), .B(n4859), .CI(
        \sub_1_root_sub_52_S2_2/carry[1] ), .CO(
        \sub_1_root_sub_52_S2_2/carry[2] ), .S(N186) );
  DFFRX1 \current_state_reg[1]  ( .D(next_state[1]), .CK(clk), .RN(n6074), 
        .QN(n5977) );
  ADDFXL \add_0_root_add_0_root_add_92_2/U1_3  ( .A(N241), .B(N235), .CI(
        \add_0_root_add_0_root_add_92_2/carry[3] ), .CO(
        \add_0_root_add_0_root_add_92_2/carry[4] ), .S(N247) );
  EDFFX1 \stringNum_reg[4]  ( .D(stringCounter[4]), .E(n3297), .CK(clk), .Q(
        n6293), .QN(\sub_1_root_add_0_root_add_92_2/n1 ) );
  ADDHXL U3788 ( .A(N170), .B(\add_0_root_add_51/carry[4] ), .CO(
        \add_0_root_add_51/carry[5] ), .S(N176) );
  ADDHXL U3786 ( .A(N169), .B(\add_0_root_add_51/carry[3] ), .CO(
        \add_0_root_add_51/carry[4] ), .S(N175) );
  ADDHXL U3784 ( .A(N167), .B(N166), .CO(\add_0_root_add_51/carry[2] ), .S(
        N173) );
  ADDHXL U3785 ( .A(N168), .B(\add_0_root_add_51/carry[2] ), .CO(
        \add_0_root_add_51/carry[3] ), .S(N174) );
  EDFFX1 \stringNum_reg[3]  ( .D(stringCounter[3]), .E(n3297), .CK(clk), .Q(
        stringNum[3]) );
  EDFFX1 \stringNum_reg[0]  ( .D(stringCounter[0]), .E(n3297), .CK(clk), .QN(
        \sub_1_root_add_0_root_add_92_2/n3 ) );
  DFFRX1 \patternCounter_reg[3]  ( .D(n1446), .CK(clk), .RN(n6421), .Q(
        patternCounter[3]), .QN(n6021) );
  ADDFXL U4682 ( .A(n4003), .B(special_locate[2]), .CI(\add_653_S2/carry[2] ), 
        .CO(\add_653_S2/carry[3] ), .S(N851) );
  ADDFXL \r685/U2_2  ( .A(stringNum[2]), .B(n4860), .CI(\r685/carry[2] ), .CO(
        \r685/carry[3] ), .S(N168) );
  ADDFXL \r685/U2_3  ( .A(stringNum[3]), .B(n6021), .CI(\r685/carry[3] ), .CO(
        \r685/carry[4] ), .S(N169) );
  ADDFXL \r685/U2_1  ( .A(stringNum[1]), .B(n4834), .CI(
        \sub_1_root_add_0_root_add_92_2/carry[1] ), .CO(\r685/carry[2] ), .S(
        N167) );
  DFFRX1 \pattern_reg[0]  ( .D(n1445), .CK(clk), .RN(n6416), .Q(pattern[0]) );
  DFFRX1 \pattern_reg[7]  ( .D(n1438), .CK(clk), .RN(n6417), .Q(pattern[7]) );
  DFFRHQX1 valid_reg ( .D(n4457), .CK(clk), .RN(n6438), .Q(n6478) );
  DFFRX1 \current_state_reg[2]  ( .D(next_state[2]), .CK(clk), .RN(n6074), .Q(
        n4848), .QN(n374) );
  DFFRHQX1 match_reg ( .D(N842), .CK(clk), .RN(n6075), .Q(n6275) );
  DFFRX1 \stringCounter_reg[3]  ( .D(n1711), .CK(clk), .RN(n6075), .Q(
        stringCounter[3]), .QN(n4853) );
  DFFRX1 \stringCounter_reg[2]  ( .D(n1713), .CK(clk), .RN(n6074), .Q(
        stringCounter[2]), .QN(n4854) );
  DFFRX1 \stringCounter_reg[0]  ( .D(n1717), .CK(clk), .RN(n6075), .Q(
        stringCounter[0]), .QN(n4856) );
  DFFSRX1 \special_locate_reg[2]  ( .D(n1722), .CK(clk), .SN(1'b1), .RN(n6075), 
        .Q(special_locate[2]), .QN(n4858) );
  DFFSRX1 \match_index_reg[2]  ( .D(n1377), .CK(clk), .SN(1'b1), .RN(n6075), 
        .Q(n4003), .QN(n452) );
  DFFSRX1 \match_index_reg[1]  ( .D(n1379), .CK(clk), .SN(1'b1), .RN(n6074), 
        .Q(n4004), .QN(n453) );
  DFFSRXL \match_index_reg[3]  ( .D(n1375), .CK(clk), .SN(1'b1), .RN(n6075), 
        .Q(n4002), .QN(n451) );
  DFFSRXL \stringCounter_reg[4]  ( .D(n1709), .CK(clk), .SN(1'b1), .RN(n6074), 
        .Q(stringCounter[4]), .QN(n4851) );
  DFFSRXL \stringCounter_reg[5]  ( .D(n1719), .CK(clk), .SN(1'b1), .RN(n6074), 
        .Q(stringCounter[5]), .QN(n4850) );
  DFFSRXL \stringData_reg[191]  ( .D(n1516), .CK(clk), .SN(1'b1), .RN(n6075), 
        .QN(n4780) );
  DFFSRXL \stringData_reg[190]  ( .D(n1517), .CK(clk), .SN(1'b1), .RN(n6074), 
        .QN(n4781) );
  DFFSRXL \stringData_reg[189]  ( .D(n1518), .CK(clk), .SN(1'b1), .RN(n6075), 
        .QN(n4782) );
  DFFSRXL \stringData_reg[188]  ( .D(n1519), .CK(clk), .SN(1'b1), .RN(n6074), 
        .QN(n4783) );
  DFFSRXL \stringData_reg[187]  ( .D(n1520), .CK(clk), .SN(1'b1), .RN(n6075), 
        .QN(n4784) );
  DFFSRXL \stringData_reg[186]  ( .D(n1521), .CK(clk), .SN(1'b1), .RN(n6074), 
        .QN(n4785) );
  DFFSRXL \stringData_reg[185]  ( .D(n1522), .CK(clk), .SN(1'b1), .RN(n6075), 
        .QN(n4786) );
  DFFSRXL \stringData_reg[184]  ( .D(n1523), .CK(clk), .SN(1'b1), .RN(n6074), 
        .QN(n4787) );
  DFFSRXL \stringData_reg[183]  ( .D(n1524), .CK(clk), .SN(1'b1), .RN(n6075), 
        .Q(stringData[183]), .QN(n4788) );
  DFFSRXL \stringData_reg[182]  ( .D(n1525), .CK(clk), .SN(1'b1), .RN(n6074), 
        .Q(stringData[182]), .QN(n4789) );
  DFFSRXL \stringData_reg[181]  ( .D(n1526), .CK(clk), .SN(1'b1), .RN(n6075), 
        .Q(stringData[181]), .QN(n4790) );
  DFFSRXL \stringData_reg[180]  ( .D(n1527), .CK(clk), .SN(1'b1), .RN(n6074), 
        .Q(stringData[180]), .QN(n4791) );
  DFFSRXL \stringData_reg[179]  ( .D(n1528), .CK(clk), .SN(1'b1), .RN(n6075), 
        .Q(stringData[179]), .QN(n4792) );
  DFFSRXL \stringData_reg[178]  ( .D(n1529), .CK(clk), .SN(1'b1), .RN(n6074), 
        .Q(stringData[178]), .QN(n4793) );
  DFFSRXL \stringData_reg[176]  ( .D(n1531), .CK(clk), .SN(1'b1), .RN(n6075), 
        .Q(stringData[176]), .QN(n4795) );
  DFFSRXL \stringData_reg[87]  ( .D(n1620), .CK(clk), .SN(1'b1), .RN(n6074), 
        .QN(n4700) );
  DFFSRXL \stringData_reg[86]  ( .D(n1621), .CK(clk), .SN(1'b1), .RN(n6075), 
        .Q(stringData[86]), .QN(n4701) );
  DFFSRXL \stringData_reg[85]  ( .D(n1622), .CK(clk), .SN(1'b1), .RN(n6074), 
        .Q(stringData[85]), .QN(n4702) );
  DFFSRXL \stringData_reg[84]  ( .D(n1623), .CK(clk), .SN(1'b1), .RN(n6075), 
        .Q(stringData[84]), .QN(n4703) );
  DFFSRXL \stringData_reg[83]  ( .D(n1624), .CK(clk), .SN(1'b1), .RN(n6074), 
        .Q(stringData[83]), .QN(n4704) );
  DFFSRXL \stringData_reg[82]  ( .D(n1625), .CK(clk), .SN(1'b1), .RN(n6075), 
        .Q(stringData[82]), .QN(n4705) );
  DFFSRXL \stringData_reg[80]  ( .D(n1627), .CK(clk), .SN(1'b1), .RN(n6074), 
        .Q(stringData[80]), .QN(n4707) );
  DFFSRXL \stringData_reg[175]  ( .D(n1532), .CK(clk), .SN(1'b1), .RN(n6075), 
        .QN(n4740) );
  DFFSRXL \stringData_reg[174]  ( .D(n1533), .CK(clk), .SN(1'b1), .RN(n6074), 
        .QN(n4741) );
  DFFSRXL \stringData_reg[173]  ( .D(n1534), .CK(clk), .SN(1'b1), .RN(n6075), 
        .QN(n4742) );
  DFFSRXL \stringData_reg[172]  ( .D(n1535), .CK(clk), .SN(1'b1), .RN(n6074), 
        .QN(n4743) );
  DFFSRXL \stringData_reg[171]  ( .D(n1536), .CK(clk), .SN(1'b1), .RN(n6075), 
        .QN(n4744) );
  DFFSRXL \stringData_reg[170]  ( .D(n1537), .CK(clk), .SN(1'b1), .RN(n6074), 
        .QN(n4745) );
  DFFSRXL \stringData_reg[168]  ( .D(n1539), .CK(clk), .SN(1'b1), .RN(n6075), 
        .QN(n4747) );
  DFFSRXL \stringData_reg[167]  ( .D(n1540), .CK(clk), .SN(1'b1), .RN(n6074), 
        .Q(stringData[167]), .QN(n4748) );
  DFFSRXL \stringData_reg[166]  ( .D(n1541), .CK(clk), .SN(1'b1), .RN(n6075), 
        .Q(stringData[166]), .QN(n4749) );
  DFFSRXL \stringData_reg[165]  ( .D(n1542), .CK(clk), .SN(1'b1), .RN(n6074), 
        .Q(stringData[165]), .QN(n4750) );
  DFFSRXL \stringData_reg[164]  ( .D(n1543), .CK(clk), .SN(1'b1), .RN(n6075), 
        .Q(stringData[164]), .QN(n4751) );
  DFFSRXL \stringData_reg[163]  ( .D(n1544), .CK(clk), .SN(1'b1), .RN(n6074), 
        .Q(stringData[163]), .QN(n4752) );
  DFFSRXL \stringData_reg[162]  ( .D(n1545), .CK(clk), .SN(1'b1), .RN(n6075), 
        .Q(stringData[162]), .QN(n4753) );
  DFFSRXL \stringData_reg[160]  ( .D(n1547), .CK(clk), .SN(1'b1), .RN(n6074), 
        .Q(stringData[160]), .QN(n4755) );
  DFFSRXL \stringData_reg[95]  ( .D(n1612), .CK(clk), .SN(1'b1), .RN(n6075), 
        .Q(stringData[95]), .QN(n4692) );
  DFFSRXL \stringData_reg[94]  ( .D(n1613), .CK(clk), .SN(1'b1), .RN(n6074), 
        .Q(stringData[94]), .QN(n4693) );
  DFFSRXL \stringData_reg[93]  ( .D(n1614), .CK(clk), .SN(1'b1), .RN(n6075), 
        .Q(stringData[93]), .QN(n4694) );
  DFFSRXL \stringData_reg[92]  ( .D(n1615), .CK(clk), .SN(1'b1), .RN(n6074), 
        .Q(stringData[92]), .QN(n4695) );
  DFFSRXL \stringData_reg[91]  ( .D(n1616), .CK(clk), .SN(1'b1), .RN(n6075), 
        .Q(stringData[91]), .QN(n4696) );
  DFFSRXL \stringData_reg[90]  ( .D(n1617), .CK(clk), .SN(1'b1), .RN(n6074), 
        .Q(stringData[90]), .QN(n4697) );
  DFFSRXL \stringData_reg[88]  ( .D(n1619), .CK(clk), .SN(1'b1), .RN(n6075), 
        .Q(stringData[88]), .QN(n4699) );
  DFFSRXL \stringData_reg[79]  ( .D(n1628), .CK(clk), .SN(1'b1), .RN(n6074), 
        .QN(n4660) );
  DFFSRXL \stringData_reg[78]  ( .D(n1629), .CK(clk), .SN(1'b1), .RN(n6075), 
        .QN(n4661) );
  DFFSRXL \stringData_reg[77]  ( .D(n1630), .CK(clk), .SN(1'b1), .RN(n6074), 
        .QN(n4662) );
  DFFSRXL \stringData_reg[76]  ( .D(n1631), .CK(clk), .SN(1'b1), .RN(n6075), 
        .QN(n4663) );
  DFFSRXL \stringData_reg[75]  ( .D(n1632), .CK(clk), .SN(1'b1), .RN(n6074), 
        .QN(n4664) );
  DFFSRXL \stringData_reg[74]  ( .D(n1633), .CK(clk), .SN(1'b1), .RN(n6075), 
        .QN(n4665) );
  DFFSRXL \stringData_reg[72]  ( .D(n1635), .CK(clk), .SN(1'b1), .RN(n6074), 
        .QN(n4667) );
  DFFSRXL \stringData_reg[71]  ( .D(n1636), .CK(clk), .SN(1'b1), .RN(n6075), 
        .QN(n4668) );
  DFFSRXL \stringData_reg[70]  ( .D(n1637), .CK(clk), .SN(1'b1), .RN(n6074), 
        .QN(n4669) );
  DFFSRXL \stringData_reg[69]  ( .D(n1638), .CK(clk), .SN(1'b1), .RN(n6075), 
        .QN(n4670) );
  DFFSRXL \stringData_reg[68]  ( .D(n1639), .CK(clk), .SN(1'b1), .RN(n6074), 
        .QN(n4671) );
  DFFSRXL \stringData_reg[67]  ( .D(n1640), .CK(clk), .SN(1'b1), .RN(n6075), 
        .QN(n4672) );
  DFFSRXL \stringData_reg[66]  ( .D(n1641), .CK(clk), .SN(1'b1), .RN(n6074), 
        .QN(n4673) );
  DFFSRXL \stringData_reg[64]  ( .D(n1643), .CK(clk), .SN(1'b1), .RN(n6075), 
        .QN(n4675) );
  DFFSRXL \stringData_reg[177]  ( .D(n1530), .CK(clk), .SN(1'b1), .RN(n6074), 
        .Q(stringData[177]), .QN(n4794) );
  DFFSRXL \stringData_reg[81]  ( .D(n1626), .CK(clk), .SN(1'b1), .RN(n6075), 
        .Q(stringData[81]), .QN(n4706) );
  DFFSRXL \stringData_reg[169]  ( .D(n1538), .CK(clk), .SN(1'b1), .RN(n6074), 
        .QN(n4746) );
  DFFSRXL \stringData_reg[161]  ( .D(n1546), .CK(clk), .SN(1'b1), .RN(n6075), 
        .Q(stringData[161]), .QN(n4754) );
  DFFSRXL \stringData_reg[89]  ( .D(n1618), .CK(clk), .SN(1'b1), .RN(n6074), 
        .Q(stringData[89]), .QN(n4698) );
  DFFSRXL \stringData_reg[73]  ( .D(n1634), .CK(clk), .SN(1'b1), .RN(n6075), 
        .QN(n4666) );
  DFFSRXL \stringData_reg[65]  ( .D(n1642), .CK(clk), .SN(1'b1), .RN(n6074), 
        .QN(n4674) );
  DFFSRXL \pattern_reg[24]  ( .D(n1421), .CK(clk), .SN(1'b1), .RN(n6075), .Q(
        pattern[24]), .QN(n4871) );
  DFFSRXL \pattern_reg[29]  ( .D(n1416), .CK(clk), .SN(1'b1), .RN(n6074), .Q(
        pattern[29]), .QN(n4867) );
  DFFSRXL \pattern_reg[27]  ( .D(n1418), .CK(clk), .SN(1'b1), .RN(n6075), .Q(
        pattern[27]), .QN(n4868) );
  DFFSRXL \pattern_reg[26]  ( .D(n1419), .CK(clk), .SN(1'b1), .RN(n6074), .Q(
        pattern[26]), .QN(n4869) );
  DFFSRXL \pattern_reg[25]  ( .D(n1420), .CK(clk), .SN(1'b1), .RN(n6075), .Q(
        pattern[25]), .QN(n4870) );
  DFFSRXL \pattern_reg[31]  ( .D(n1414), .CK(clk), .SN(1'b1), .RN(n6074), .Q(
        pattern[31]) );
  DFFSRXL \pattern_reg[30]  ( .D(n1415), .CK(clk), .SN(1'b1), .RN(n6075), .Q(
        pattern[30]) );
  DFFSRXL \pattern_reg[28]  ( .D(n1417), .CK(clk), .SN(1'b1), .RN(n6074), .Q(
        pattern[28]) );
  DFFSRXL \pattern_reg[23]  ( .D(n1422), .CK(clk), .SN(1'b1), .RN(n6075), .Q(
        pattern[23]), .QN(n4872) );
  DFFSRXL \pattern_reg[22]  ( .D(n1423), .CK(clk), .SN(1'b1), .RN(n6074), .Q(
        pattern[22]), .QN(n4873) );
  DFFSRXL \pattern_reg[20]  ( .D(n1425), .CK(clk), .SN(1'b1), .RN(n6075), .Q(
        pattern[20]), .QN(n4874) );
  DFFSRXL \pattern_reg[16]  ( .D(n1429), .CK(clk), .SN(1'b1), .RN(n6074), .QN(
        n4555) );
  DFFSRXL \pattern_reg[21]  ( .D(n1424), .CK(clk), .SN(1'b1), .RN(n6075), .Q(
        pattern[21]), .QN(n4875) );
  DFFSRXL \pattern_reg[19]  ( .D(n1426), .CK(clk), .SN(1'b1), .RN(n6074), .Q(
        pattern[19]), .QN(n4876) );
  DFFSRXL \pattern_reg[18]  ( .D(n1427), .CK(clk), .SN(1'b1), .RN(n6075), .Q(
        pattern[18]), .QN(n4877) );
  DFFSRXL \pattern_reg[17]  ( .D(n1428), .CK(clk), .SN(1'b1), .RN(n6074), .Q(
        pattern[17]), .QN(n4878) );
  DFFSRXL \stringData_reg[7]  ( .D(n1700), .CK(clk), .SN(1'b1), .RN(n6075), 
        .QN(n4684) );
  DFFSRXL \stringData_reg[6]  ( .D(n1701), .CK(clk), .SN(1'b1), .RN(n6074), 
        .QN(n4685) );
  DFFSRXL \stringData_reg[4]  ( .D(n1703), .CK(clk), .SN(1'b1), .RN(n6075), 
        .QN(n4686) );
  DFFSRXL \stringData_reg[2]  ( .D(n1705), .CK(clk), .SN(1'b1), .RN(n6074), 
        .QN(n4688) );
  DFFSRXL \stringData_reg[0]  ( .D(n1707), .CK(clk), .SN(1'b1), .RN(n6075), 
        .QN(n4690) );
  DFFSRXL \stringData_reg[3]  ( .D(n1704), .CK(clk), .SN(1'b1), .RN(n6074), 
        .QN(n4687) );
  DFFSRXL \stringData_reg[1]  ( .D(n1706), .CK(clk), .SN(1'b1), .RN(n6075), 
        .QN(n4689) );
  DFFSRXL \stringData_reg[5]  ( .D(n1702), .CK(clk), .SN(1'b1), .RN(n6074), 
        .Q(stringData[5]) );
  DFFSRXL \stringData_reg[231]  ( .D(n1476), .CK(clk), .SN(1'b1), .RN(n6075), 
        .QN(n4820) );
  DFFSRXL \stringData_reg[230]  ( .D(n1477), .CK(clk), .SN(1'b1), .RN(n6074), 
        .QN(n4821) );
  DFFSRXL \stringData_reg[229]  ( .D(n1478), .CK(clk), .SN(1'b1), .RN(n6075), 
        .QN(n4822) );
  DFFSRXL \stringData_reg[228]  ( .D(n1479), .CK(clk), .SN(1'b1), .RN(n6074), 
        .QN(n4823) );
  DFFSRXL \stringData_reg[227]  ( .D(n1480), .CK(clk), .SN(1'b1), .RN(n6075), 
        .QN(n4824) );
  DFFSRXL \stringData_reg[226]  ( .D(n1481), .CK(clk), .SN(1'b1), .RN(n6074), 
        .QN(n4825) );
  DFFSRXL \stringData_reg[225]  ( .D(n1482), .CK(clk), .SN(1'b1), .RN(n6075), 
        .QN(n4826) );
  DFFSRXL \stringData_reg[224]  ( .D(n1483), .CK(clk), .SN(1'b1), .RN(n6074), 
        .QN(n4827) );
  DFFSRXL \stringData_reg[223]  ( .D(n1484), .CK(clk), .SN(1'b1), .RN(n6075), 
        .QN(n4764) );
  DFFSRXL \stringData_reg[222]  ( .D(n1485), .CK(clk), .SN(1'b1), .RN(n6074), 
        .QN(n4765) );
  DFFSRXL \stringData_reg[221]  ( .D(n1486), .CK(clk), .SN(1'b1), .RN(n6075), 
        .QN(n4766) );
  DFFSRXL \stringData_reg[220]  ( .D(n1487), .CK(clk), .SN(1'b1), .RN(n6074), 
        .QN(n4767) );
  DFFSRXL \stringData_reg[219]  ( .D(n1488), .CK(clk), .SN(1'b1), .RN(n6075), 
        .QN(n4768) );
  DFFSRXL \stringData_reg[218]  ( .D(n1489), .CK(clk), .SN(1'b1), .RN(n6074), 
        .QN(n4769) );
  DFFSRXL \stringData_reg[217]  ( .D(n1490), .CK(clk), .SN(1'b1), .RN(n6075), 
        .QN(n4770) );
  DFFSRXL \stringData_reg[216]  ( .D(n1491), .CK(clk), .SN(1'b1), .RN(n6074), 
        .QN(n4771) );
  DFFSRXL \stringData_reg[215]  ( .D(n1492), .CK(clk), .SN(1'b1), .RN(n6075), 
        .Q(stringData[215]), .QN(n4772) );
  DFFSRXL \stringData_reg[214]  ( .D(n1493), .CK(clk), .SN(1'b1), .RN(n6074), 
        .QN(n4773) );
  DFFSRXL \stringData_reg[213]  ( .D(n1494), .CK(clk), .SN(1'b1), .RN(n6075), 
        .QN(n4774) );
  DFFSRXL \stringData_reg[212]  ( .D(n1495), .CK(clk), .SN(1'b1), .RN(n6074), 
        .QN(n4775) );
  DFFSRXL \stringData_reg[211]  ( .D(n1496), .CK(clk), .SN(1'b1), .RN(n6075), 
        .QN(n4776) );
  DFFSRXL \stringData_reg[210]  ( .D(n1497), .CK(clk), .SN(1'b1), .RN(n6074), 
        .QN(n4777) );
  DFFSRXL \stringData_reg[209]  ( .D(n1498), .CK(clk), .SN(1'b1), .RN(n6075), 
        .QN(n4778) );
  DFFSRXL \stringData_reg[208]  ( .D(n1499), .CK(clk), .SN(1'b1), .RN(n6074), 
        .QN(n4779) );
  DFFSRXL \stringData_reg[207]  ( .D(n1500), .CK(clk), .SN(1'b1), .RN(n6075), 
        .Q(stringData[207]), .QN(n4724) );
  DFFSRXL \stringData_reg[206]  ( .D(n1501), .CK(clk), .SN(1'b1), .RN(n6074), 
        .Q(stringData[206]), .QN(n4725) );
  DFFSRXL \stringData_reg[204]  ( .D(n1503), .CK(clk), .SN(1'b1), .RN(n6075), 
        .Q(stringData[204]), .QN(n4727) );
  DFFSRXL \stringData_reg[203]  ( .D(n1504), .CK(clk), .SN(1'b1), .RN(n6074), 
        .Q(stringData[203]), .QN(n4728) );
  DFFSRXL \stringData_reg[202]  ( .D(n1505), .CK(clk), .SN(1'b1), .RN(n6075), 
        .Q(stringData[202]), .QN(n4729) );
  DFFSRXL \stringData_reg[201]  ( .D(n1506), .CK(clk), .SN(1'b1), .RN(n6074), 
        .Q(stringData[201]), .QN(n4730) );
  DFFSRXL \stringData_reg[200]  ( .D(n1507), .CK(clk), .SN(1'b1), .RN(n6075), 
        .Q(stringData[200]), .QN(n4731) );
  DFFSRXL \stringData_reg[197]  ( .D(n1510), .CK(clk), .SN(1'b1), .RN(n6074), 
        .QN(n4734) );
  DFFSRXL \stringData_reg[195]  ( .D(n1512), .CK(clk), .SN(1'b1), .RN(n6075), 
        .QN(n4736) );
  DFFSRXL \stringData_reg[193]  ( .D(n1514), .CK(clk), .SN(1'b1), .RN(n6074), 
        .QN(n4738) );
  DFFSRXL \stringData_reg[239]  ( .D(n1468), .CK(clk), .SN(1'b1), .RN(n6075), 
        .Q(stringData[239]), .QN(n4812) );
  DFFSRXL \stringData_reg[238]  ( .D(n1469), .CK(clk), .SN(1'b1), .RN(n6074), 
        .Q(stringData[238]), .QN(n4813) );
  DFFSRXL \stringData_reg[237]  ( .D(n1470), .CK(clk), .SN(1'b1), .RN(n6075), 
        .Q(stringData[237]), .QN(n4814) );
  DFFSRXL \stringData_reg[236]  ( .D(n1471), .CK(clk), .SN(1'b1), .RN(n6074), 
        .Q(stringData[236]), .QN(n4815) );
  DFFSRXL \stringData_reg[235]  ( .D(n1472), .CK(clk), .SN(1'b1), .RN(n6075), 
        .Q(stringData[235]), .QN(n4816) );
  DFFSRXL \stringData_reg[234]  ( .D(n1473), .CK(clk), .SN(1'b1), .RN(n6074), 
        .Q(stringData[234]), .QN(n4817) );
  DFFSRXL \stringData_reg[232]  ( .D(n1475), .CK(clk), .SN(1'b1), .RN(n6075), 
        .Q(stringData[232]), .QN(n4819) );
  DFFSRXL \stringData_reg[63]  ( .D(n1644), .CK(clk), .SN(1'b1), .RN(n6074), 
        .QN(n4708) );
  DFFSRXL \stringData_reg[62]  ( .D(n1645), .CK(clk), .SN(1'b1), .RN(n6075), 
        .QN(n4709) );
  DFFSRXL \stringData_reg[61]  ( .D(n1646), .CK(clk), .SN(1'b1), .RN(n6074), 
        .QN(n4710) );
  DFFSRXL \stringData_reg[60]  ( .D(n1647), .CK(clk), .SN(1'b1), .RN(n6075), 
        .QN(n4711) );
  DFFSRXL \stringData_reg[59]  ( .D(n1648), .CK(clk), .SN(1'b1), .RN(n6074), 
        .QN(n4712) );
  DFFSRXL \stringData_reg[58]  ( .D(n1649), .CK(clk), .SN(1'b1), .RN(n6075), 
        .QN(n4713) );
  DFFSRXL \stringData_reg[56]  ( .D(n1651), .CK(clk), .SN(1'b1), .RN(n6074), 
        .QN(n4715) );
  DFFSRXL \stringData_reg[47]  ( .D(n1660), .CK(clk), .SN(1'b1), .RN(n6075), 
        .QN(n4676) );
  DFFSRXL \stringData_reg[46]  ( .D(n1661), .CK(clk), .SN(1'b1), .RN(n6074), 
        .QN(n4677) );
  DFFSRXL \stringData_reg[45]  ( .D(n1662), .CK(clk), .SN(1'b1), .RN(n6075), 
        .QN(n4678) );
  DFFSRXL \stringData_reg[44]  ( .D(n1663), .CK(clk), .SN(1'b1), .RN(n6074), 
        .QN(n4679) );
  DFFSRXL \stringData_reg[43]  ( .D(n1664), .CK(clk), .SN(1'b1), .RN(n6075), 
        .QN(n4680) );
  DFFSRXL \stringData_reg[42]  ( .D(n1665), .CK(clk), .SN(1'b1), .RN(n6074), 
        .QN(n4681) );
  DFFSRXL \stringData_reg[40]  ( .D(n1667), .CK(clk), .SN(1'b1), .RN(n6075), 
        .QN(n4683) );
  DFFSRXL \stringData_reg[233]  ( .D(n1474), .CK(clk), .SN(1'b1), .RN(n6074), 
        .Q(stringData[233]), .QN(n4818) );
  DFFSRXL \stringData_reg[41]  ( .D(n1666), .CK(clk), .SN(1'b1), .RN(n6075), 
        .QN(n4682) );
  DFFSRXL \stringData_reg[205]  ( .D(n1502), .CK(clk), .SN(1'b1), .RN(n6074), 
        .Q(stringData[205]), .QN(n4726) );
  DFFSRXL \stringData_reg[199]  ( .D(n1508), .CK(clk), .SN(1'b1), .RN(n6075), 
        .QN(n4732) );
  DFFSRXL \stringData_reg[198]  ( .D(n1509), .CK(clk), .SN(1'b1), .RN(n6074), 
        .QN(n4733) );
  DFFSRXL \stringData_reg[196]  ( .D(n1511), .CK(clk), .SN(1'b1), .RN(n6075), 
        .QN(n4735) );
  DFFSRXL \stringData_reg[194]  ( .D(n1513), .CK(clk), .SN(1'b1), .RN(n6074), 
        .QN(n4737) );
  DFFSRXL \stringData_reg[192]  ( .D(n1515), .CK(clk), .SN(1'b1), .RN(n6075), 
        .QN(n4739) );
  DFFSRXL \stringData_reg[159]  ( .D(n1548), .CK(clk), .SN(1'b1), .RN(n6074), 
        .QN(n4796) );
  DFFSRXL \stringData_reg[158]  ( .D(n1549), .CK(clk), .SN(1'b1), .RN(n6075), 
        .QN(n4797) );
  DFFSRXL \stringData_reg[157]  ( .D(n1550), .CK(clk), .SN(1'b1), .RN(n6074), 
        .QN(n4798) );
  DFFSRXL \stringData_reg[156]  ( .D(n1551), .CK(clk), .SN(1'b1), .RN(n6075), 
        .QN(n4799) );
  DFFSRXL \stringData_reg[155]  ( .D(n1552), .CK(clk), .SN(1'b1), .RN(n6074), 
        .QN(n4800) );
  DFFSRXL \stringData_reg[154]  ( .D(n1553), .CK(clk), .SN(1'b1), .RN(n6075), 
        .QN(n4801) );
  DFFSRXL \stringData_reg[152]  ( .D(n1555), .CK(clk), .SN(1'b1), .RN(n6074), 
        .QN(n4803) );
  DFFSRXL \stringData_reg[151]  ( .D(n1556), .CK(clk), .SN(1'b1), .RN(n6075), 
        .Q(stringData[151]), .QN(n4804) );
  DFFSRXL \stringData_reg[150]  ( .D(n1557), .CK(clk), .SN(1'b1), .RN(n6074), 
        .Q(stringData[150]), .QN(n4805) );
  DFFSRXL \stringData_reg[149]  ( .D(n1558), .CK(clk), .SN(1'b1), .RN(n6075), 
        .Q(stringData[149]), .QN(n4806) );
  DFFSRXL \stringData_reg[148]  ( .D(n1559), .CK(clk), .SN(1'b1), .RN(n6074), 
        .Q(stringData[148]), .QN(n4807) );
  DFFSRXL \stringData_reg[147]  ( .D(n1560), .CK(clk), .SN(1'b1), .RN(n6075), 
        .Q(stringData[147]), .QN(n4808) );
  DFFSRXL \stringData_reg[146]  ( .D(n1561), .CK(clk), .SN(1'b1), .RN(n6074), 
        .Q(stringData[146]), .QN(n4809) );
  DFFSRXL \stringData_reg[144]  ( .D(n1563), .CK(clk), .SN(1'b1), .RN(n6075), 
        .Q(stringData[144]), .QN(n4811) );
  DFFSRXL \stringData_reg[135]  ( .D(n1572), .CK(clk), .SN(1'b1), .RN(n6074), 
        .QN(n4756) );
  DFFSRXL \stringData_reg[134]  ( .D(n1573), .CK(clk), .SN(1'b1), .RN(n6075), 
        .QN(n4757) );
  DFFSRXL \stringData_reg[133]  ( .D(n1574), .CK(clk), .SN(1'b1), .RN(n6074), 
        .Q(stringData[133]), .QN(n4758) );
  DFFSRXL \stringData_reg[132]  ( .D(n1575), .CK(clk), .SN(1'b1), .RN(n6075), 
        .QN(n4759) );
  DFFSRXL \stringData_reg[131]  ( .D(n1576), .CK(clk), .SN(1'b1), .RN(n6074), 
        .QN(n4760) );
  DFFSRXL \stringData_reg[130]  ( .D(n1577), .CK(clk), .SN(1'b1), .RN(n6075), 
        .QN(n4761) );
  DFFSRXL \stringData_reg[128]  ( .D(n1579), .CK(clk), .SN(1'b1), .RN(n6074), 
        .QN(n4763) );
  DFFSRXL \stringData_reg[111]  ( .D(n1596), .CK(clk), .SN(1'b1), .RN(n6075), 
        .Q(stringData[111]), .QN(n4652) );
  DFFSRXL \stringData_reg[110]  ( .D(n1597), .CK(clk), .SN(1'b1), .RN(n6074), 
        .Q(stringData[110]), .QN(n4653) );
  DFFSRXL \stringData_reg[109]  ( .D(n1598), .CK(clk), .SN(1'b1), .RN(n6075), 
        .Q(stringData[109]), .QN(n4654) );
  DFFSRXL \stringData_reg[108]  ( .D(n1599), .CK(clk), .SN(1'b1), .RN(n6074), 
        .Q(stringData[108]), .QN(n4655) );
  DFFSRXL \stringData_reg[107]  ( .D(n1600), .CK(clk), .SN(1'b1), .RN(n6075), 
        .Q(stringData[107]), .QN(n4656) );
  DFFSRXL \stringData_reg[106]  ( .D(n1601), .CK(clk), .SN(1'b1), .RN(n6074), 
        .Q(stringData[106]), .QN(n4657) );
  DFFSRXL \stringData_reg[104]  ( .D(n1603), .CK(clk), .SN(1'b1), .RN(n6075), 
        .Q(stringData[104]), .QN(n4659) );
  DFFSRXL \stringData_reg[55]  ( .D(n1652), .CK(clk), .SN(1'b1), .RN(n6074), 
        .QN(n4716) );
  DFFSRXL \stringData_reg[54]  ( .D(n1653), .CK(clk), .SN(1'b1), .RN(n6075), 
        .QN(n4717) );
  DFFSRXL \stringData_reg[53]  ( .D(n1654), .CK(clk), .SN(1'b1), .RN(n6074), 
        .QN(n4718) );
  DFFSRXL \stringData_reg[52]  ( .D(n1655), .CK(clk), .SN(1'b1), .RN(n6075), 
        .QN(n4719) );
  DFFSRXL \stringData_reg[51]  ( .D(n1656), .CK(clk), .SN(1'b1), .RN(n6074), 
        .QN(n4720) );
  DFFSRXL \stringData_reg[50]  ( .D(n1657), .CK(clk), .SN(1'b1), .RN(n6075), 
        .QN(n4721) );
  DFFSRXL \stringData_reg[48]  ( .D(n1659), .CK(clk), .SN(1'b1), .RN(n6074), 
        .QN(n4723) );
  DFFSRXL \stringData_reg[153]  ( .D(n1554), .CK(clk), .SN(1'b1), .RN(n6075), 
        .QN(n4802) );
  DFFSRXL \stringData_reg[145]  ( .D(n1562), .CK(clk), .SN(1'b1), .RN(n6074), 
        .Q(stringData[145]), .QN(n4810) );
  DFFRX2 \patternCounter_reg[1]  ( .D(n1448), .CK(clk), .RN(n6074), .Q(
        patternCounter[1]), .QN(n4834) );
  DFFSRX2 \special_locate_reg[1]  ( .D(n1450), .CK(clk), .SN(1'b1), .RN(n6074), 
        .Q(special_locate[1]), .QN(n4859) );
  DFFSRX1 special_reg ( .D(n1449), .CK(clk), .SN(1'b1), .RN(n6074), .Q(special), .QN(n4857) );
  DFFSRX1 \stringCounter_reg[1]  ( .D(n1715), .CK(clk), .SN(1'b1), .RN(n6075), 
        .Q(stringCounter[1]), .QN(n4855) );
  DFFRX2 \patternCounter_reg[2]  ( .D(n1447), .CK(clk), .RN(n6075), .Q(
        patternCounter[2]), .QN(n4860) );
  DFFRX1 \match_index_reg[4]  ( .D(n1720), .CK(clk), .RN(n6427), .Q(n6288), 
        .QN(n449) );
  DFFSRX1 \patternCounter_reg[0]  ( .D(n1723), .CK(clk), .SN(1'b1), .RN(n6075), 
        .Q(patternCounter[0]), .QN(n6004) );
  OAI221X1 U4790 ( .A0(n5017), .A1(n4684), .B0(n6457), .B1(n5717), .C0(n5718), 
        .Y(n5353) );
  NAND3BX2 U4791 ( .AN(n5039), .B(n5038), .C(n6006), .Y(n5037) );
  NOR2X6 U4792 ( .A(n4458), .B(n4857), .Y(n6006) );
  OAI221X4 U4793 ( .A0(n4632), .A1(n5404), .B0(n4633), .B1(n5403), .C0(n6027), 
        .Y(n5361) );
  INVX2 U4794 ( .A(n5362), .Y(n4633) );
  AOI222XL U4795 ( .A0(n6305), .A1(n4797), .B0(n6306), .B1(n4765), .C0(n6307), 
        .C1(n4693), .Y(n5804) );
  OAI222XL U4796 ( .A0(n5619), .A1(n6383), .B0(n5620), .B1(n6381), .C0(n6465), 
        .C1(n5621), .Y(n5586) );
  OAI222XL U4797 ( .A0(n5627), .A1(n6383), .B0(n5529), .B1(n6381), .C0(n6465), 
        .C1(n5530), .Y(n5573) );
  OAI222XL U4798 ( .A0(n5623), .A1(n6383), .B0(n5561), .B1(n6381), .C0(n6465), 
        .C1(n5562), .Y(n5582) );
  OAI222XL U4799 ( .A0(n5620), .A1(n6387), .B0(n5619), .B1(n6385), .C0(
        match_index[1]), .C1(n4616), .Y(n5647) );
  OAI222XL U4800 ( .A0(n5616), .A1(n6387), .B0(n5615), .B1(n6385), .C0(
        match_index[1]), .C1(n4611), .Y(n5650) );
  OAI222XL U4801 ( .A0(n5529), .A1(n6387), .B0(n5627), .B1(n6385), .C0(
        match_index[1]), .C1(n4643), .Y(n5658) );
  OAI222XL U4802 ( .A0(n5844), .A1(n6387), .B0(n5787), .B1(n6386), .C0(
        match_index[1]), .C1(n4613), .Y(n5827) );
  OAI222XL U4803 ( .A0(n5783), .A1(n6383), .B0(n5545), .B1(n6382), .C0(n6464), 
        .C1(n5546), .Y(n5635) );
  OAI22XL U4804 ( .A0(n6456), .A1(n5827), .B0(n6297), .B1(n5786), .Y(n5321) );
  OAI222XL U4805 ( .A0(n5615), .A1(n6383), .B0(n5616), .B1(n6381), .C0(n6465), 
        .C1(n5617), .Y(n5590) );
  OAI222XL U4806 ( .A0(n4585), .A1(n5370), .B0(n4876), .B1(n5371), .C0(n5374), 
        .C1(n5372), .Y(n5335) );
  BUFX4 U4807 ( .A(n5655), .Y(n6370) );
  OAI221XL U4808 ( .A0(n4608), .A1(n5404), .B0(n4610), .B1(n5403), .C0(n6028), 
        .Y(n5350) );
  OAI221XL U4809 ( .A0(n5017), .A1(n4690), .B0(n6457), .B1(n5720), .C0(n5721), 
        .Y(n5362) );
  OAI222XL U4810 ( .A0(n6384), .A1(n5587), .B0(n5588), .B1(n6382), .C0(n6465), 
        .C1(n5589), .Y(n5522) );
  AO22X1 U4811 ( .A0(n6297), .A1(n5725), .B0(n5726), .B1(n6458), .Y(n5357) );
  OAI211X1 U4812 ( .A0(n5384), .A1(n5979), .B0(n5683), .C0(n5684), .Y(n5442)
         );
  CLKINVX1 U4813 ( .A(n5732), .Y(n4612) );
  NOR3BX1 U4814 ( .AN(n4932), .B(n4853), .C(stringCounter[2]), .Y(n4939) );
  NOR3BX1 U4815 ( .AN(n4954), .B(n4854), .C(stringCounter[3]), .Y(n4956) );
  CLKINVX4 U4816 ( .A(n4993), .Y(n4465) );
  CLKBUFX3 U4817 ( .A(n6466), .Y(n6471) );
  NAND2X2 U4818 ( .A(n4465), .B(chardata[4]), .Y(n4983) );
  NAND2X2 U4819 ( .A(n4465), .B(chardata[6]), .Y(n4985) );
  NAND2X2 U4820 ( .A(n4465), .B(chardata[7]), .Y(n4986) );
  NAND2X2 U4821 ( .A(n4465), .B(chardata[3]), .Y(n4982) );
  NAND2X2 U4822 ( .A(n4465), .B(chardata[1]), .Y(n4979) );
  NAND2X2 U4823 ( .A(n4465), .B(chardata[0]), .Y(n4978) );
  NAND2X2 U4824 ( .A(n4465), .B(chardata[5]), .Y(n4984) );
  NAND2X2 U4825 ( .A(n4465), .B(chardata[2]), .Y(n4981) );
  INVX1 U4826 ( .A(n5001), .Y(n4458) );
  AOI222XL U4827 ( .A0(n4847), .A1(n4845), .B0(n5068), .B1(n4848), .C0(n5069), 
        .C1(n4849), .Y(n5063) );
  INVX3 U4828 ( .A(n6313), .Y(n4449) );
  OAI2BB2XL U4829 ( .B0(n6299), .B1(n5032), .A0N(pattern_after[54]), .A1N(
        n6299), .Y(n1330) );
  OAI22XL U4830 ( .A0(n6067), .A1(n5024), .B0(n6299), .B1(n5030), .Y(n1344) );
  OAI22XL U4831 ( .A0(n6299), .A1(n5033), .B0(n6066), .B1(n5024), .Y(n1323) );
  OAI22XL U4832 ( .A0(n6005), .A1(n5024), .B0(n6299), .B1(n5029), .Y(n1351) );
  OAI22XL U4833 ( .A0(n6060), .A1(n5024), .B0(n6299), .B1(n5027), .Y(n1365) );
  OAI22XL U4834 ( .A0(n6068), .A1(n5024), .B0(n6299), .B1(n5031), .Y(n1337) );
  OAI22XL U4835 ( .A0(n6069), .A1(n5024), .B0(n6299), .B1(n5028), .Y(n1353) );
  OAI22XL U4836 ( .A0(n6052), .A1(n5024), .B0(n6299), .B1(n5018), .Y(n1367) );
  INVX1 U4837 ( .A(n5382), .Y(n4639) );
  OAI222X2 U4838 ( .A0(n5619), .A1(n6381), .B0(n5757), .B1(n6383), .C0(n6465), 
        .C1(n4616), .Y(n5717) );
  INVX3 U4839 ( .A(n6370), .Y(n6380) );
  AND2X2 U4840 ( .A(n451), .B(n6288), .Y(n6292) );
  INVX1 U4841 ( .A(n6370), .Y(n6379) );
  NAND2X4 U4842 ( .A(n6477), .B(n6349), .Y(n5655) );
  INVXL U4843 ( .A(n5036), .Y(n4544) );
  BUFX4 U4844 ( .A(n449), .Y(n6349) );
  NAND3X2 U4845 ( .A(n5065), .B(n4468), .C(n374), .Y(n5064) );
  NAND2XL U4846 ( .A(patternCounter[2]), .B(n4858), .Y(n5090) );
  NOR2XL U4847 ( .A(n4859), .B(n4858), .Y(N241) );
  NOR3XL U4848 ( .A(patternCounter[2]), .B(patternCounter[3]), .C(n4834), .Y(
        n5153) );
  INVXL U4849 ( .A(n6275), .Y(n6071) );
  INVX12 U4850 ( .A(n6071), .Y(match) );
  INVX3 U4851 ( .A(n4836), .Y(n6073) );
  INVX16 U4852 ( .A(n6073), .Y(n6074) );
  INVX16 U4853 ( .A(n6073), .Y(n6075) );
  BUFX12 U5052 ( .A(n6478), .Y(valid) );
  CLKBUFX3 U5053 ( .A(n4454), .Y(n6300) );
  CLKINVX1 U5054 ( .A(n5019), .Y(n4454) );
  NOR3BX2 U5055 ( .AN(n6287), .B(n5127), .C(n5330), .Y(n5315) );
  CLKBUFX3 U5056 ( .A(n4460), .Y(n6298) );
  CLKINVX1 U5057 ( .A(n4999), .Y(n4460) );
  CLKINVX1 U5058 ( .A(n5364), .Y(n4619) );
  CLKBUFX3 U5059 ( .A(n5702), .Y(n6360) );
  INVX3 U5060 ( .A(n6354), .Y(n6352) );
  OAI221X4 U5061 ( .A0(n5017), .A1(n4685), .B0(n6457), .B1(n5705), .C0(n5706), 
        .Y(n5351) );
  AOI222XL U5062 ( .A0(n5698), .A1(n5699), .B0(n4641), .B1(n5700), .C0(n4642), 
        .C1(n5701), .Y(n5697) );
  AOI222XL U5063 ( .A0(n5698), .A1(n5722), .B0(n4634), .B1(n5700), .C0(n4635), 
        .C1(n5701), .Y(n5721) );
  CLKINVX1 U5064 ( .A(n5807), .Y(n4631) );
  CLKBUFX3 U5065 ( .A(next_state[0]), .Y(n6276) );
  INVX3 U5066 ( .A(n5026), .Y(n4456) );
  CLKINVX1 U5067 ( .A(n5351), .Y(n4610) );
  NOR2X1 U5068 ( .A(match_index[1]), .B(n4642), .Y(n6283) );
  OAI22XL U5069 ( .A0(n4610), .A1(n5417), .B0(n5983), .B1(n5418), .Y(n5419) );
  INVXL U5070 ( .A(n6380), .Y(n6277) );
  NAND2X2 U5071 ( .A(n6291), .B(n6308), .Y(n5024) );
  OR3X2 U5072 ( .A(n6281), .B(n6282), .C(n6283), .Y(n5674) );
  NAND2X1 U5073 ( .A(n6288), .B(n4002), .Y(n5656) );
  CLKINVX1 U5074 ( .A(n5037), .Y(n6289) );
  OAI22XL U5075 ( .A0(n6458), .A1(n5674), .B0(n6295), .B1(n5696), .Y(n5382) );
  NAND2BX1 U5076 ( .AN(n4976), .B(n4465), .Y(n4997) );
  AND2XL U5077 ( .A(pattern[7]), .B(n4615), .Y(n6286) );
  AND2X1 U5078 ( .A(n5698), .B(n5707), .Y(n6278) );
  AND2X2 U5079 ( .A(n4630), .B(n5700), .Y(n6279) );
  AND2XL U5080 ( .A(n4631), .B(n5701), .Y(n6280) );
  NOR3X1 U5081 ( .A(n6278), .B(n6279), .C(n6280), .Y(n5706) );
  CLKINVX1 U5082 ( .A(n5024), .Y(n4455) );
  NOR2X2 U5083 ( .A(n6381), .B(match_index[0]), .Y(n5700) );
  NAND3X1 U5084 ( .A(n6289), .B(n6290), .C(n5036), .Y(n6291) );
  CLKBUFX3 U5085 ( .A(n6357), .Y(n6362) );
  OAI222XL U5086 ( .A0(n6387), .A1(n5648), .B0(n4637), .B1(n6386), .C0(
        match_index[1]), .C1(n4638), .Y(n5672) );
  OAI222XL U5087 ( .A0(n6361), .A1(n4671), .B0(n6369), .B1(n4735), .C0(n6352), 
        .C1(n4759), .Y(n5699) );
  CLKBUFX3 U5088 ( .A(n4970), .Y(n6308) );
  NAND4X1 U5089 ( .A(n5408), .B(n5409), .C(n5410), .D(n5411), .Y(n5125) );
  CLKINVX1 U5090 ( .A(n5355), .Y(n4640) );
  NOR2X1 U5091 ( .A(n6388), .B(n5581), .Y(n6281) );
  NOR2X1 U5092 ( .A(n4641), .B(n6385), .Y(n6282) );
  INVX1 U5093 ( .A(n5752), .Y(n4642) );
  NOR2X2 U5094 ( .A(n6383), .B(match_index[0]), .Y(n5698) );
  INVXL U5095 ( .A(n5102), .Y(n4518) );
  NAND2X1 U5096 ( .A(n6464), .B(n6472), .Y(n5574) );
  CLKBUFX3 U5097 ( .A(n6467), .Y(n6472) );
  OAI21X4 U5098 ( .A0(n375), .A1(isstring), .B0(n5066), .Y(n5065) );
  CLKBUFX3 U5099 ( .A(n453), .Y(n6461) );
  AND2XL U5100 ( .A(pattern[0]), .B(n4633), .Y(n6284) );
  AND2X2 U5101 ( .A(n5422), .B(n5417), .Y(n6285) );
  NOR3X1 U5102 ( .A(n6284), .B(n6285), .C(n6286), .Y(n5410) );
  CLKINVX1 U5103 ( .A(n5353), .Y(n4615) );
  INVX1 U5104 ( .A(n5429), .Y(n4471) );
  NAND2X1 U5105 ( .A(n5001), .B(n4971), .Y(n4993) );
  BUFX8 U5106 ( .A(n452), .Y(n6469) );
  NOR3BX4 U5107 ( .AN(next_state[0]), .B(next_state[1]), .C(next_state[2]), 
        .Y(n5001) );
  INVX3 U5108 ( .A(n6373), .Y(n6372) );
  INVX3 U5109 ( .A(n6374), .Y(n6371) );
  INVX3 U5110 ( .A(n6309), .Y(n4450) );
  INVX3 U5111 ( .A(n6312), .Y(n4453) );
  INVX3 U5112 ( .A(n6310), .Y(n4451) );
  INVX3 U5113 ( .A(n6311), .Y(n4452) );
  CLKINVX1 U5114 ( .A(n5240), .Y(n4585) );
  INVX3 U5115 ( .A(n4980), .Y(n4464) );
  INVX3 U5116 ( .A(n6315), .Y(n4463) );
  NOR3X1 U5117 ( .A(n5311), .B(n5312), .C(n5126), .Y(n5303) );
  OAI22X1 U5118 ( .A0(n6455), .A1(n5647), .B0(n6297), .B1(n5672), .Y(n5323) );
  INVX3 U5119 ( .A(n6292), .Y(n6351) );
  INVX3 U5120 ( .A(n5000), .Y(n4459) );
  INVX3 U5121 ( .A(n4996), .Y(n4462) );
  INVX3 U5122 ( .A(n4998), .Y(n4461) );
  CLKINVX1 U5123 ( .A(n5360), .Y(n4617) );
  CLKINVX1 U5124 ( .A(n5035), .Y(n6290) );
  CLKBUFX3 U5125 ( .A(n5656), .Y(n6367) );
  OAI32X1 U5126 ( .A0(n5133), .A1(n5131), .A2(n5086), .B0(n4648), .B1(n5134), 
        .Y(n5077) );
  OAI22X1 U5127 ( .A0(n6455), .A1(n5653), .B0(n6297), .B1(n5670), .Y(n5242) );
  OAI22X1 U5128 ( .A0(n6455), .A1(n5650), .B0(n6295), .B1(n5673), .Y(n5333) );
  INVX3 U5129 ( .A(n6354), .Y(n6353) );
  OAI22XL U5130 ( .A0(n5096), .A1(n4976), .B0(n5097), .B1(n5075), .Y(n5095) );
  OAI211X1 U5131 ( .A0(n5094), .A1(n5095), .B0(n4468), .C0(n4847), .Y(n5011)
         );
  OAI211X1 U5132 ( .A0(n4507), .A1(n4995), .B0(n5139), .C0(n5140), .Y(n5094)
         );
  OAI22XL U5133 ( .A0(n4640), .A1(n5417), .B0(n6010), .B1(n5418), .Y(n5416) );
  NOR3X1 U5134 ( .A(n5406), .B(n5125), .C(n5407), .Y(n5397) );
  NOR3X1 U5135 ( .A(n5287), .B(n5086), .C(n5288), .Y(n5279) );
  NOR3X1 U5136 ( .A(n5299), .B(n5085), .C(n5300), .Y(n5291) );
  NOR3X1 U5137 ( .A(n5275), .B(n5084), .C(n5276), .Y(n5266) );
  CLKINVX1 U5138 ( .A(n4918), .Y(n4426) );
  AOI222XL U5139 ( .A0(n5698), .A1(n5711), .B0(n4626), .B1(n5700), .C0(n4625), 
        .C1(n5701), .Y(n5710) );
  AOI222XL U5140 ( .A0(n5698), .A1(n5715), .B0(n4627), .B1(n5700), .C0(n4624), 
        .C1(n5701), .Y(n5714) );
  OAI222X1 U5141 ( .A0(n6388), .A1(n5585), .B0(n4634), .B1(n6386), .C0(
        match_index[1]), .C1(n4635), .Y(n5670) );
  OAI221XL U5142 ( .A0(n6008), .A1(n5418), .B0(n5417), .B1(n5357), .C0(n5012), 
        .Y(n5423) );
  AOI222XL U5143 ( .A0(n5698), .A1(n5719), .B0(n5700), .B1(n4637), .C0(n5701), 
        .C1(n4638), .Y(n5718) );
  OAI22XL U5144 ( .A0(n4612), .A1(n5417), .B0(n6031), .B1(n5418), .Y(n5424) );
  OAI22XL U5145 ( .A0(n4619), .A1(n5417), .B0(n6015), .B1(n5418), .Y(n5420) );
  OAI22XL U5146 ( .A0(n4617), .A1(n5417), .B0(n6016), .B1(n5418), .Y(n5421) );
  OA22X1 U5147 ( .A0(n6457), .A1(n5786), .B0(n6297), .B1(n5733), .Y(n5375) );
  OAI221XL U5148 ( .A0(n5017), .A1(n4688), .B0(n6457), .B1(n5733), .C0(n5734), 
        .Y(n5732) );
  CLKINVX1 U5149 ( .A(n5443), .Y(n4475) );
  OAI222XL U5150 ( .A0(n5430), .A1(n5431), .B0(n5432), .B1(n5433), .C0(n5434), 
        .C1(n5435), .Y(n5429) );
  NAND2X1 U5151 ( .A(n6349), .B(n4002), .Y(n5702) );
  OAI32X1 U5152 ( .A0(n5099), .A1(patternCounter[2]), .A2(patternCounter[1]), 
        .B0(n5100), .B1(n4976), .Y(n5098) );
  AOI221XL U5153 ( .A0(n4830), .A1(n4556), .B0(n4832), .B1(n4553), .C0(n5098), 
        .Y(n5097) );
  OAI221X1 U5154 ( .A0(n6353), .A1(n4791), .B0(n6372), .B1(n4719), .C0(n5754), 
        .Y(n5575) );
  NAND4X1 U5155 ( .A(n5603), .B(n5604), .C(n5605), .D(n5606), .Y(n5449) );
  NAND4X1 U5156 ( .A(n5637), .B(n5638), .C(n5639), .D(n5640), .Y(n5448) );
  NAND2XL U5157 ( .A(n6359), .B(match_index[2]), .Y(n5577) );
  CLKINVX1 U5158 ( .A(n5525), .Y(n6390) );
  CLKINVX1 U5159 ( .A(n5525), .Y(n6389) );
  CLKBUFX2 U5160 ( .A(n6357), .Y(n6361) );
  NAND2X1 U5161 ( .A(n6472), .B(match_index[1]), .Y(n5528) );
  NAND2XL U5162 ( .A(match_index[2]), .B(match_index[1]), .Y(n5525) );
  NOR2XL U5163 ( .A(n5655), .B(n6471), .Y(n5580) );
  XNOR2X1 U5164 ( .A(n5333), .B(n5334), .Y(n6287) );
  OAI32XL U5165 ( .A0(n5137), .A1(n5131), .A2(n5084), .B0(n4648), .B1(n5138), 
        .Y(n5078) );
  OAI22XL U5166 ( .A0(n6456), .A1(n5843), .B0(n6296), .B1(n5827), .Y(n5840) );
  OAI22XL U5167 ( .A0(n6458), .A1(n5819), .B0(n6295), .B1(n5782), .Y(n5325) );
  OAI22XL U5168 ( .A0(n6455), .A1(n5618), .B0(n6295), .B1(n5647), .Y(n5644) );
  OAI22XL U5169 ( .A0(n6455), .A1(n5614), .B0(n6295), .B1(n5650), .Y(n5642) );
  OAI22XL U5170 ( .A0(n6455), .A1(n5626), .B0(n6296), .B1(n5658), .Y(n5645) );
  XNOR2XL U5171 ( .A(n5358), .B(n4612), .Y(n5141) );
  CLKINVX3 U5172 ( .A(n4994), .Y(n4466) );
  CLKBUFX2 U5173 ( .A(n6363), .Y(n6369) );
  XOR2XL U5174 ( .A(n5327), .B(n5328), .Y(n5317) );
  XOR2XL U5175 ( .A(n5325), .B(n5326), .Y(n5318) );
  XOR2XL U5176 ( .A(n5321), .B(n5322), .Y(n5320) );
  XNOR2XL U5177 ( .A(n5374), .B(n5335), .Y(n5366) );
  XNOR2XL U5178 ( .A(n5381), .B(n5326), .Y(n5380) );
  XNOR2XL U5179 ( .A(n5369), .B(n5328), .Y(n5368) );
  XOR2XL U5180 ( .A(n5323), .B(n5324), .Y(n5319) );
  XOR2XL U5181 ( .A(n5360), .B(n5712), .Y(n5689) );
  XOR2XL U5182 ( .A(n5364), .B(n5708), .Y(n5690) );
  XOR2XL U5183 ( .A(n5351), .B(n5704), .Y(n5691) );
  CLKINVX3 U5184 ( .A(n6314), .Y(n4467) );
  CLKBUFX2 U5185 ( .A(n6363), .Y(n6368) );
  NAND2XL U5186 ( .A(n6464), .B(match_index[2]), .Y(n5576) );
  INVX16 U5187 ( .A(n6463), .Y(match_index[1]) );
  OAI22XL U5188 ( .A0(n6022), .A1(n5635), .B0(n6297), .B1(n5636), .Y(n5632) );
  OAI22XL U5189 ( .A0(n6022), .A1(n5590), .B0(n6295), .B1(n5614), .Y(n5610) );
  OAI22XL U5190 ( .A0(n6022), .A1(n5582), .B0(n6296), .B1(n5622), .Y(n5612) );
  OAI22XL U5191 ( .A0(n6022), .A1(n5586), .B0(n6296), .B1(n5618), .Y(n5608) );
  OAI22XL U5192 ( .A0(n6022), .A1(n5573), .B0(n6297), .B1(n5626), .Y(n5611) );
  CLKINVX1 U5193 ( .A(n6453), .Y(n6294) );
  NAND2XL U5194 ( .A(n6354), .B(match_index[2]), .Y(n5578) );
  OAI22XL U5195 ( .A0(n6456), .A1(n5540), .B0(n6295), .B1(n5870), .Y(n5884) );
  OAI22XL U5196 ( .A0(n6022), .A1(n5522), .B0(n6297), .B1(n5586), .Y(n5571) );
  OAI22XL U5197 ( .A0(n6022), .A1(n5558), .B0(n6297), .B1(n5582), .Y(n5568) );
  OAI22XL U5198 ( .A0(n6455), .A1(n5523), .B0(match_index[0]), .B1(n5573), .Y(
        n5570) );
  XOR2XL U5199 ( .A(n6472), .B(n5393), .Y(n5390) );
  OAI32XL U5200 ( .A0(n5345), .A1(n5127), .A2(n5131), .B0(n4648), .B1(n5236), 
        .Y(n5344) );
  NAND2XL U5201 ( .A(n6295), .B(n6464), .Y(n5927) );
  XOR2X1 U5202 ( .A(n5040), .B(n5041), .Y(n5036) );
  XNOR2XL U5203 ( .A(n5381), .B(n5356), .Y(n5407) );
  NOR4XL U5204 ( .A(n5105), .B(n5106), .C(n5102), .D(n5107), .Y(n5104) );
  OAI222XL U5205 ( .A0(n6387), .A1(n5814), .B0(n4627), .B1(n6386), .C0(
        match_index[1]), .C1(n4624), .Y(n5778) );
  OAI222XL U5206 ( .A0(n5820), .A1(n6387), .B0(n4629), .B1(n6386), .C0(
        match_index[1]), .C1(n4621), .Y(n5782) );
  OAI222XL U5207 ( .A0(n6388), .A1(n5775), .B0(n4626), .B1(n6386), .C0(
        match_index[1]), .C1(n4625), .Y(n5682) );
  OAI222XL U5208 ( .A0(n6387), .A1(n5828), .B0(n4628), .B1(n6386), .C0(
        match_index[1]), .C1(n4623), .Y(n5786) );
  OAI221XL U5209 ( .A0(n4614), .A1(n5404), .B0(n4615), .B1(n5403), .C0(n6029), 
        .Y(n5352) );
  OAI221XL U5210 ( .A0(n4639), .A1(n5404), .B0(n4640), .B1(n5403), .C0(n6030), 
        .Y(n5354) );
  OAI22X1 U5211 ( .A0(n6458), .A1(n5673), .B0(n6296), .B1(n5705), .Y(n5384) );
  OAI22XL U5212 ( .A0(n6458), .A1(n5672), .B0(n6297), .B1(n5717), .Y(n5383) );
  OAI22X1 U5213 ( .A0(n6458), .A1(n5670), .B0(n6297), .B1(n5720), .Y(n5373) );
  NAND3XL U5214 ( .A(n4860), .B(n6021), .C(n4465), .Y(n4988) );
  AOI211XL U5215 ( .A0(n4527), .A1(n4547), .B0(n5083), .C0(n4518), .Y(n5081)
         );
  INVXL U5216 ( .A(n5086), .Y(n4527) );
  OAI222XL U5217 ( .A0(n5381), .A1(n5372), .B0(n4577), .B1(n5370), .C0(n4554), 
        .C1(n4875), .Y(n5326) );
  OAI222XL U5218 ( .A0(n4581), .A1(n5370), .B0(n4878), .B1(n5371), .C0(n5369), 
        .C1(n5372), .Y(n5328) );
  OAI222XL U5219 ( .A0(n4594), .A1(n5370), .B0(n4877), .B1(n5371), .C0(n5375), 
        .C1(n5372), .Y(n5322) );
  OAI222XL U5220 ( .A0(n5858), .A1(n6387), .B0(n5772), .B1(n6386), .C0(
        match_index[1]), .C1(n4620), .Y(n5681) );
  OAI222XL U5221 ( .A0(n5545), .A1(n6387), .B0(n5783), .B1(n6386), .C0(
        match_index[1]), .C1(n4622), .Y(n5819) );
  OAI221XL U5222 ( .A0(n4561), .A1(n5370), .B0(n4632), .B1(n5372), .C0(n4555), 
        .Y(n5336) );
  OAI221XL U5223 ( .A0(n4587), .A1(n5370), .B0(n4614), .B1(n5372), .C0(n4872), 
        .Y(n5324) );
  OAI221XL U5224 ( .A0(n4567), .A1(n5370), .B0(n4639), .B1(n5372), .C0(n4874), 
        .Y(n5332) );
  OAI221XL U5225 ( .A0(n4597), .A1(n5370), .B0(n4608), .B1(n5372), .C0(n4873), 
        .Y(n5334) );
  OAI2BB1XL U5226 ( .A0N(n5045), .A1N(n4511), .B0(n5014), .Y(n5044) );
  NOR2X1 U5227 ( .A(n5017), .B(n5012), .Y(n5149) );
  NOR3BX1 U5228 ( .AN(n4954), .B(n4853), .C(n4854), .Y(n4966) );
  NOR3BX1 U5229 ( .AN(n4932), .B(n4853), .C(n4854), .Y(n4944) );
  XNOR2XL U5230 ( .A(n5356), .B(n5357), .Y(n5148) );
  OAI32XL U5231 ( .A0(n5444), .A1(n5442), .A2(n5462), .B0(n5463), .B1(n4551), 
        .Y(n5459) );
  XOR2XL U5232 ( .A(n5242), .B(n5243), .Y(n5224) );
  XOR2XL U5233 ( .A(n5240), .B(n5241), .Y(n5225) );
  XOR2XL U5234 ( .A(n5355), .B(n5693), .Y(n5692) );
  XOR2XL U5235 ( .A(n6464), .B(N245), .Y(n5049) );
  XOR2XL U5236 ( .A(n5239), .B(n4597), .Y(n5235) );
  XOR2XL U5237 ( .A(n5238), .B(n4567), .Y(n5237) );
  XOR2XL U5238 ( .A(n5240), .B(n5812), .Y(n5676) );
  XOR2XL U5239 ( .A(n5327), .B(n5678), .Y(n5677) );
  OR2X1 U5240 ( .A(n4971), .B(n4458), .Y(n4912) );
  NAND4XL U5241 ( .A(n4582), .B(n4580), .C(n5440), .D(n5496), .Y(n5431) );
  NAND2XL U5242 ( .A(next_state[1]), .B(n6276), .Y(n4970) );
  AOI2BB2XL U5243 ( .B0(n6390), .B1(n5602), .A0N(n6384), .A1N(n4626), .Y(n5878) );
  OAI222XL U5244 ( .A0(n5779), .A1(n6383), .B0(n5850), .B1(n6382), .C0(n6461), 
        .C1(n5886), .Y(n5870) );
  OAI222XL U5245 ( .A0(n5772), .A1(n6383), .B0(n5858), .B1(n6382), .C0(n6463), 
        .C1(n5882), .Y(n5599) );
  OAI221XL U5246 ( .A0(n5591), .A1(n6385), .B0(n6382), .B1(n5651), .C0(n5652), 
        .Y(n5614) );
  AOI2BB2XL U5247 ( .B0(n6389), .B1(n5593), .A0N(n6384), .A1N(n4630), .Y(n5652) );
  OAI221XL U5248 ( .A0(n5587), .A1(n6385), .B0(n6382), .B1(n5648), .C0(n5649), 
        .Y(n5618) );
  OA22XL U5249 ( .A0(n6384), .A1(n4637), .B0(n6388), .B1(n5588), .Y(n5649) );
  OAI221XL U5250 ( .A0(n5575), .A1(n6385), .B0(n6382), .B1(n5581), .C0(n5659), 
        .Y(n5626) );
  AOI2BB2XL U5251 ( .B0(n6389), .B1(n5508), .A0N(n6384), .A1N(n4641), .Y(n5659) );
  OAI221XL U5252 ( .A0(n5583), .A1(n6385), .B0(n6382), .B1(n5585), .C0(n5654), 
        .Y(n5622) );
  AOI2BB2XL U5253 ( .B0(n6389), .B1(n5503), .A0N(n6384), .A1N(n4634), .Y(n5654) );
  OAI221XL U5254 ( .A0(n5830), .A1(n6385), .B0(n6382), .B1(n5828), .C0(n5865), 
        .Y(n5843) );
  AOI2BB2XL U5255 ( .B0(n6390), .B1(n5866), .A0N(n6384), .A1N(n4628), .Y(n5865) );
  OAI221XL U5256 ( .A0(n6047), .A1(n5298), .B0(n4574), .B1(n5297), .C0(n5130), 
        .Y(n5244) );
  NAND2X1 U5257 ( .A(n5012), .B(n5417), .Y(n5418) );
  OAI32XL U5258 ( .A0(n5466), .A1(n5445), .A2(n5056), .B0(n5448), .B1(n5467), 
        .Y(n5465) );
  XOR2XL U5259 ( .A(n5233), .B(n4587), .Y(n5230) );
  OAI221XL U5260 ( .A0(n5816), .A1(n6385), .B0(n6382), .B1(n5814), .C0(n5871), 
        .Y(n5849) );
  AOI2BB2XL U5261 ( .B0(n6389), .B1(n5872), .A0N(n6384), .A1N(n4627), .Y(n5871) );
  OAI221XL U5262 ( .A0(n5822), .A1(n6385), .B0(n6382), .B1(n5820), .C0(n5837), 
        .Y(n5636) );
  AOI2BB2XL U5263 ( .B0(n6390), .B1(n5513), .A0N(n6384), .A1N(n4629), .Y(n5837) );
  OAI222XL U5264 ( .A0(n6384), .A1(n5591), .B0(n4607), .B1(n6381), .C0(n6465), 
        .C1(n5592), .Y(n5531) );
  OAI222XL U5265 ( .A0(n6384), .A1(n5583), .B0(n4601), .B1(n6381), .C0(n6465), 
        .C1(n5501), .Y(n5558) );
  OAI222XL U5266 ( .A0(n6384), .A1(n5575), .B0(n4602), .B1(n6382), .C0(n453), 
        .C1(n5507), .Y(n5523) );
  OAI222XL U5267 ( .A0(n6384), .A1(n5830), .B0(n4606), .B1(n6382), .C0(n6465), 
        .C1(n5894), .Y(n5548) );
  OAI222XL U5268 ( .A0(n6384), .A1(n5816), .B0(n4605), .B1(n6382), .C0(n6461), 
        .C1(n5888), .Y(n5540) );
  OAI222XL U5269 ( .A0(n5787), .A1(n6383), .B0(n5844), .B1(n6382), .C0(n6461), 
        .C1(n5892), .Y(n5864) );
  OAI221XL U5270 ( .A0(n6048), .A1(n5285), .B0(n4573), .B1(n5286), .C0(n5133), 
        .Y(n5253) );
  INVXL U5271 ( .A(n5445), .Y(n4537) );
  OAI222XL U5272 ( .A0(n6384), .A1(n5600), .B0(n4604), .B1(n6381), .C0(n6465), 
        .C1(n5601), .Y(n5555) );
  OAI221XL U5273 ( .A0(n6056), .A1(n5273), .B0(n4578), .B1(n5274), .C0(n5137), 
        .Y(n5184) );
  OAI22XL U5274 ( .A0(n6455), .A1(n5499), .B0(n6296), .B1(n5558), .Y(n5342) );
  OAI22XL U5275 ( .A0(match_index[0]), .A1(n5523), .B0(n6456), .B1(n5505), .Y(
        n5518) );
  OAI22XL U5276 ( .A0(match_index[0]), .A1(n5531), .B0(n6456), .B1(n5532), .Y(
        n5262) );
  NAND2X1 U5277 ( .A(n5695), .B(n5724), .Y(n5694) );
  INVXL U5278 ( .A(n5125), .Y(n4609) );
  AOI222X1 U5279 ( .A0(N168), .A1(n4515), .B0(N187), .B1(n4512), .C0(N174), 
        .C1(n5484), .Y(n5393) );
  AOI222X1 U5280 ( .A0(N167), .A1(n4515), .B0(N186), .B1(n4512), .C0(N173), 
        .C1(n5484), .Y(n5452) );
  CLKBUFX3 U5281 ( .A(n4843), .Y(n6394) );
  CLKBUFX3 U5282 ( .A(n4844), .Y(n6392) );
  CLKBUFX3 U5283 ( .A(n4842), .Y(n6396) );
  CLKBUFX3 U5284 ( .A(n4841), .Y(n6398) );
  CLKBUFX3 U5285 ( .A(n4840), .Y(n6400) );
  CLKBUFX3 U5286 ( .A(n4839), .Y(n6402) );
  CLKBUFX3 U5287 ( .A(n4838), .Y(n6404) );
  CLKBUFX3 U5288 ( .A(n4837), .Y(n6406) );
  XOR2XL U5289 ( .A(match_index[2]), .B(N246), .Y(n5054) );
  AO21XL U5290 ( .A0(n6359), .A1(\add_653_S2/carry[3] ), .B0(n6356), .Y(n4919)
         );
  NOR2X2 U5291 ( .A(n4855), .B(n4856), .Y(n4931) );
  AOI22XL U5292 ( .A0(n6358), .A1(stringData[114]), .B0(stringData[242]), .B1(
        n6365), .Y(n5895) );
  AOI22XL U5293 ( .A0(n6358), .A1(stringData[115]), .B0(stringData[243]), .B1(
        n6365), .Y(n5889) );
  INVXL U5294 ( .A(n5043), .Y(n4470) );
  AOI33XL U5295 ( .A0(n5047), .A1(n4468), .A2(n374), .B0(n4511), .B1(n5045), 
        .B2(n5014), .Y(n5046) );
  OAI221XL U5296 ( .A0(n6353), .A1(n4783), .B0(n6372), .B1(n4711), .C0(n5749), 
        .Y(n5629) );
  AOI22XL U5297 ( .A0(n6359), .A1(stringData[124]), .B0(stringData[252]), .B1(
        n6364), .Y(n5749) );
  OAI221XL U5298 ( .A0(n6353), .A1(n4781), .B0(n6372), .B1(n4709), .C0(n5956), 
        .Y(n5803) );
  AOI22XL U5299 ( .A0(n6358), .A1(stringData[126]), .B0(stringData[254]), .B1(
        n6364), .Y(n5956) );
  OAI221XL U5300 ( .A0(n6352), .A1(n4787), .B0(n6372), .B1(n4715), .C0(n5793), 
        .Y(n5625) );
  AOI22XL U5301 ( .A0(n6358), .A1(stringData[121]), .B0(stringData[249]), .B1(
        n6365), .Y(n5912) );
  AOI22XL U5302 ( .A0(n6358), .A1(stringData[123]), .B0(stringData[251]), .B1(
        n6365), .Y(n5921) );
  AOI22XL U5303 ( .A0(n6358), .A1(stringData[122]), .B0(stringData[250]), .B1(
        n6364), .Y(n5946) );
  INVXL U5304 ( .A(n5017), .Y(n4649) );
  NOR3XL U5305 ( .A(n4911), .B(n5977), .C(n6276), .Y(n5015) );
  AOI22XL U5306 ( .A0(n6358), .A1(stringData[117]), .B0(stringData[245]), .B1(
        n6365), .Y(n5903) );
  AOI22XL U5307 ( .A0(N856), .A1(n4918), .B0(N850), .B1(n4449), .Y(n5007) );
  AOI22XL U5308 ( .A0(N857), .A1(n4918), .B0(N851), .B1(n4449), .Y(n5008) );
  OAI22XL U5309 ( .A0(n6004), .A1(n4846), .B0(ispattern), .B1(n6308), .Y(n4972) );
  NOR3BX1 U5310 ( .AN(n4954), .B(n4853), .C(stringCounter[2]), .Y(n4961) );
  NOR3BX1 U5311 ( .AN(n4932), .B(n4854), .C(stringCounter[3]), .Y(n4934) );
  NOR3BX1 U5312 ( .AN(n4954), .B(stringCounter[2]), .C(stringCounter[3]), .Y(
        n4950) );
  NOR3BX1 U5313 ( .AN(n4932), .B(stringCounter[2]), .C(stringCounter[3]), .Y(
        n4925) );
  NAND2X1 U5314 ( .A(n6006), .B(chardata[7]), .Y(n5033) );
  NAND2X1 U5315 ( .A(n6006), .B(chardata[4]), .Y(n5030) );
  NAND2X1 U5316 ( .A(n6006), .B(chardata[0]), .Y(n5018) );
  NAND2X1 U5317 ( .A(n6006), .B(chardata[3]), .Y(n5029) );
  NAND2X1 U5318 ( .A(n6006), .B(chardata[1]), .Y(n5027) );
  NAND2X1 U5319 ( .A(n6006), .B(chardata[5]), .Y(n5031) );
  NAND2X1 U5320 ( .A(n6006), .B(chardata[2]), .Y(n5028) );
  NAND2X1 U5321 ( .A(n6006), .B(chardata[6]), .Y(n5032) );
  XOR2XL U5322 ( .A(n5968), .B(n5369), .Y(n5771) );
  XOR2XL U5323 ( .A(n5729), .B(n4612), .Y(n5685) );
  XOR2XL U5324 ( .A(n5357), .B(n5723), .Y(n5686) );
  AOI22XL U5325 ( .A0(n6358), .A1(stringData[125]), .B0(stringData[253]), .B1(
        n6365), .Y(n5898) );
  OAI211XL U5326 ( .A0(n6476), .A1(n4920), .B0(n5009), .C0(n5010), .Y(n1375)
         );
  NAND3XL U5327 ( .A(n4449), .B(n6476), .C(\add_653_S2/carry[3] ), .Y(n5009)
         );
  AOI2BB2XL U5328 ( .B0(N858), .B1(n4918), .A0N(n5958), .A1N(n4916), .Y(n5010)
         );
  XOR2XL U5329 ( .A(n5971), .B(n5375), .Y(n5768) );
  XOR2XL U5330 ( .A(n5969), .B(n5381), .Y(n5769) );
  XOR2XL U5331 ( .A(n5970), .B(n5374), .Y(n5770) );
  OAI221XL U5332 ( .A0(n6301), .A1(n4803), .B0(n6302), .B1(n4771), .C0(n5624), 
        .Y(n5562) );
  AOI22XL U5333 ( .A0(stringData[88]), .A1(n6303), .B0(n5625), .B1(n6473), .Y(
        n5624) );
  OAI221XL U5334 ( .A0(n6301), .A1(n4799), .B0(n6302), .B1(n4767), .C0(n5628), 
        .Y(n5530) );
  AOI22XL U5335 ( .A0(stringData[92]), .A1(n6303), .B0(n5629), .B1(n6468), .Y(
        n5628) );
  OAI221XL U5336 ( .A0(n6301), .A1(n4796), .B0(n6302), .B1(n4764), .C0(n5933), 
        .Y(n5621) );
  AOI22XL U5337 ( .A0(stringData[95]), .A1(n6303), .B0(n5759), .B1(n6474), .Y(
        n5933) );
  OAI221XL U5338 ( .A0(n6301), .A1(n4797), .B0(n6302), .B1(n4765), .C0(n5955), 
        .Y(n5617) );
  AOI22XL U5339 ( .A0(stringData[94]), .A1(n6303), .B0(n5803), .B1(n6474), .Y(
        n5955) );
  OAI221XL U5340 ( .A0(n6301), .A1(n4798), .B0(n6302), .B1(n4766), .C0(n5897), 
        .Y(n5546) );
  AOI22XL U5341 ( .A0(stringData[93]), .A1(n6303), .B0(n5835), .B1(n6474), .Y(
        n5897) );
  OAI221XL U5342 ( .A0(n6301), .A1(n4800), .B0(n6302), .B1(n4768), .C0(n5920), 
        .Y(n5886) );
  AOI22XL U5343 ( .A0(stringData[91]), .A1(n6303), .B0(n5852), .B1(n6474), .Y(
        n5920) );
  OAI221XL U5344 ( .A0(n6301), .A1(n4802), .B0(n6302), .B1(n4770), .C0(n5911), 
        .Y(n5882) );
  AOI22XL U5345 ( .A0(stringData[89]), .A1(n6303), .B0(n5860), .B1(n6468), .Y(
        n5911) );
  AOI2BB2XL U5346 ( .B0(n4774), .B1(n6288), .A0N(stringData[149]), .A1N(n6477), 
        .Y(n5902) );
  AOI2BB2XL U5347 ( .B0(n4778), .B1(n6288), .A0N(stringData[145]), .A1N(n6476), 
        .Y(n5907) );
  AOI2BB2XL U5348 ( .B0(n4775), .B1(match_index[4]), .A0N(stringData[148]), 
        .A1N(n6476), .Y(n5660) );
  AOI2BB2XL U5349 ( .B0(n4779), .B1(match_index[4]), .A0N(stringData[144]), 
        .A1N(n6476), .Y(n5657) );
  AOI2BB2XL U5350 ( .B0(n4773), .B1(n6288), .A0N(stringData[150]), .A1N(n6476), 
        .Y(n5951) );
  AOI2BB2XL U5351 ( .B0(n4777), .B1(n6288), .A0N(stringData[146]), .A1N(n6476), 
        .Y(n5941) );
  OAI221XL U5352 ( .A0(n6301), .A1(n4748), .B0(n6302), .B1(n4820), .C0(n5936), 
        .Y(n5589) );
  OAI221XL U5353 ( .A0(n6301), .A1(n4755), .B0(n6302), .B1(n4827), .C0(n5584), 
        .Y(n5501) );
  OAI221XL U5354 ( .A0(n6301), .A1(n4751), .B0(n6302), .B1(n4823), .C0(n5579), 
        .Y(n5507) );
  AOI22XL U5355 ( .A0(stringData[100]), .A1(n6303), .B0(n5581), .B1(n6472), 
        .Y(n5579) );
  OAI221XL U5356 ( .A0(n6301), .A1(n4750), .B0(n6302), .B1(n4822), .C0(n5901), 
        .Y(n5512) );
  OAI221XL U5357 ( .A0(n6301), .A1(n4752), .B0(n6302), .B1(n4824), .C0(n5917), 
        .Y(n5888) );
  OAI221XL U5358 ( .A0(n6301), .A1(n4749), .B0(n6302), .B1(n4821), .C0(n5952), 
        .Y(n5592) );
  OAI221XL U5359 ( .A0(n6301), .A1(n4753), .B0(n6302), .B1(n4825), .C0(n5942), 
        .Y(n5894) );
  OAI221XL U5360 ( .A0(n6301), .A1(n4801), .B0(n6302), .B1(n4769), .C0(n5945), 
        .Y(n5892) );
  AOI22XL U5361 ( .A0(stringData[90]), .A1(n6303), .B0(n5846), .B1(n6468), .Y(
        n5945) );
  XOR2XL U5362 ( .A(match_index[3]), .B(n5392), .Y(n5391) );
  OAI221XL U5363 ( .A0(n6301), .A1(n4754), .B0(n6302), .B1(n4826), .C0(n5908), 
        .Y(n5601) );
  OAI21XL U5364 ( .A0(n5475), .A1(n5487), .B0(n5488), .Y(n5394) );
  OAI21XL U5365 ( .A0(n5475), .A1(n5485), .B0(n5486), .Y(n5392) );
  OAI222XL U5366 ( .A0(n5471), .A1(n5472), .B0(n4516), .B1(n5473), .C0(n5474), 
        .C1(n5475), .Y(n5461) );
  OAI221XL U5367 ( .A0(n5914), .A1(n5498), .B0(n6297), .B1(n5539), .C0(n5915), 
        .Y(n5123) );
  OAI221XL U5368 ( .A0(n5905), .A1(n5498), .B0(n6297), .B1(n5554), .C0(n5906), 
        .Y(n5121) );
  OAI221XL U5369 ( .A0(n5504), .A1(n5498), .B0(n6295), .B1(n5505), .C0(n5506), 
        .Y(n5169) );
  OAI221XL U5370 ( .A0(n5497), .A1(n5498), .B0(n6297), .B1(n5499), .C0(n5500), 
        .Y(n5168) );
  OAI221XL U5371 ( .A0(n5509), .A1(n5498), .B0(n6295), .B1(n5510), .C0(n5511), 
        .Y(n5260) );
  AOI211XL U5372 ( .A0(n6376), .A1(n6007), .B0(n5930), .C0(n6365), .Y(n5929)
         );
  NAND3X1 U5373 ( .A(pattern_after[17]), .B(n5825), .C(pattern_after[19]), .Y(
        n5679) );
  CLKINVX1 U5374 ( .A(chardata[1]), .Y(n4843) );
  NAND3X1 U5375 ( .A(pattern_after[25]), .B(n5855), .C(pattern_after[27]), .Y(
        n5833) );
  NAND3X1 U5376 ( .A(pattern_after[33]), .B(n5876), .C(pattern_after[35]), .Y(
        n5634) );
  NAND3X1 U5377 ( .A(pattern_after[41]), .B(n5891), .C(pattern_after[43]), .Y(
        n5597) );
  CLKINVX1 U5378 ( .A(chardata[0]), .Y(n4844) );
  CLKINVX1 U5379 ( .A(chardata[2]), .Y(n4842) );
  CLKINVX1 U5380 ( .A(chardata[3]), .Y(n4841) );
  CLKINVX1 U5381 ( .A(chardata[4]), .Y(n4840) );
  CLKINVX1 U5382 ( .A(chardata[5]), .Y(n4839) );
  CLKINVX1 U5383 ( .A(chardata[6]), .Y(n4838) );
  CLKINVX1 U5384 ( .A(chardata[7]), .Y(n4837) );
  NAND2X1 U5385 ( .A(n374), .B(n375), .Y(n4911) );
  NOR3X1 U5386 ( .A(n4849), .B(n374), .C(n4468), .Y(n5014) );
  NAND3X1 U5387 ( .A(n4848), .B(n4849), .C(n5977), .Y(n5016) );
  NOR2X2 U5388 ( .A(n4855), .B(stringCounter[0]), .Y(n4929) );
  NOR2X2 U5389 ( .A(stringCounter[0]), .B(stringCounter[1]), .Y(n4924) );
  NOR2X2 U5390 ( .A(n4856), .B(stringCounter[1]), .Y(n4927) );
  INVX16 U5391 ( .A(n6349), .Y(match_index[4]) );
  NOR2X1 U5392 ( .A(n4550), .B(n5041), .Y(n5035) );
  INVX3 U5393 ( .A(n6363), .Y(n6364) );
  INVX3 U5394 ( .A(n6367), .Y(n6365) );
  INVX3 U5395 ( .A(n6368), .Y(n6366) );
  INVX3 U5396 ( .A(n6389), .Y(n6388) );
  INVX3 U5397 ( .A(n6390), .Y(n6387) );
  NAND2X2 U5398 ( .A(n6389), .B(n6365), .Y(n5526) );
  CLKBUFX3 U5399 ( .A(n5746), .Y(n6305) );
  NOR2X1 U5400 ( .A(n6351), .B(match_index[2]), .Y(n5746) );
  CLKBUFX3 U5401 ( .A(n5747), .Y(n6306) );
  NOR2X1 U5402 ( .A(n5656), .B(match_index[2]), .Y(n5747) );
  CLKBUFX3 U5403 ( .A(n5748), .Y(n6307) );
  NOR2X1 U5404 ( .A(n6360), .B(match_index[2]), .Y(n5748) );
  INVX3 U5405 ( .A(n6357), .Y(n6359) );
  INVX3 U5406 ( .A(n6360), .Y(n6358) );
  NAND2X2 U5407 ( .A(n6374), .B(n5698), .Y(n5017) );
  CLKBUFX3 U5408 ( .A(n5528), .Y(n6386) );
  CLKBUFX3 U5409 ( .A(n5577), .Y(n6301) );
  CLKBUFX3 U5410 ( .A(n5528), .Y(n6385) );
  CLKBUFX3 U5411 ( .A(n5578), .Y(n6302) );
  NAND2X2 U5412 ( .A(n6390), .B(n6296), .Y(n5498) );
  NAND2BX2 U5413 ( .AN(n6386), .B(n6297), .Y(n5502) );
  CLKBUFX3 U5414 ( .A(n6448), .Y(n6417) );
  CLKBUFX3 U5415 ( .A(n6447), .Y(n6418) );
  CLKBUFX3 U5416 ( .A(n6447), .Y(n6419) );
  CLKBUFX3 U5417 ( .A(n6446), .Y(n6420) );
  CLKBUFX3 U5418 ( .A(n6446), .Y(n6421) );
  CLKBUFX3 U5419 ( .A(n6445), .Y(n6422) );
  CLKBUFX3 U5420 ( .A(n6445), .Y(n6423) );
  CLKBUFX3 U5421 ( .A(n6450), .Y(n6414) );
  CLKBUFX3 U5422 ( .A(n6449), .Y(n6415) );
  CLKBUFX3 U5423 ( .A(n6448), .Y(n6416) );
  CLKBUFX3 U5424 ( .A(n6439), .Y(n6433) );
  CLKBUFX3 U5425 ( .A(n6439), .Y(n6434) );
  CLKBUFX3 U5426 ( .A(n6407), .Y(n6435) );
  CLKBUFX3 U5427 ( .A(n6449), .Y(n6436) );
  CLKBUFX3 U5428 ( .A(n6407), .Y(n6437) );
  CLKBUFX3 U5429 ( .A(n6444), .Y(n6424) );
  CLKBUFX3 U5430 ( .A(n6443), .Y(n6425) );
  CLKBUFX3 U5431 ( .A(n6443), .Y(n6426) );
  CLKBUFX3 U5432 ( .A(n6442), .Y(n6427) );
  CLKBUFX3 U5433 ( .A(n6442), .Y(n6428) );
  CLKBUFX3 U5434 ( .A(n6441), .Y(n6429) );
  CLKBUFX3 U5435 ( .A(n6441), .Y(n6430) );
  CLKBUFX3 U5436 ( .A(n6440), .Y(n6431) );
  CLKBUFX3 U5437 ( .A(n6440), .Y(n6432) );
  CLKBUFX3 U5438 ( .A(n6450), .Y(n6438) );
  CLKBUFX3 U5439 ( .A(n4455), .Y(n6299) );
  CLKBUFX3 U5440 ( .A(n5656), .Y(n6363) );
  INVX16 U5441 ( .A(n6471), .Y(match_index[2]) );
  NAND4X1 U5442 ( .A(n5346), .B(n5347), .C(n5348), .D(n5349), .Y(n5236) );
  NOR4X1 U5443 ( .A(n5377), .B(n5378), .C(n5379), .D(n5380), .Y(n5346) );
  NOR4X1 U5444 ( .A(n5365), .B(n5366), .C(n5367), .D(n5368), .Y(n5347) );
  NOR4X1 U5445 ( .A(n5151), .B(n5152), .C(n5150), .D(n5141), .Y(n5348) );
  CLKINVX1 U5446 ( .A(n5321), .Y(n4594) );
  CLKINVX1 U5447 ( .A(n5325), .Y(n4577) );
  CLKINVX1 U5448 ( .A(n5327), .Y(n4581) );
  CLKINVX1 U5449 ( .A(n5242), .Y(n4561) );
  CLKINVX1 U5450 ( .A(n5323), .Y(n4587) );
  CLKINVX1 U5451 ( .A(n5331), .Y(n4567) );
  CLKINVX1 U5452 ( .A(n5333), .Y(n4597) );
  CLKBUFX3 U5453 ( .A(n5576), .Y(n6381) );
  CLKBUFX3 U5454 ( .A(n5574), .Y(n6383) );
  CLKBUFX3 U5455 ( .A(n6380), .Y(n6374) );
  CLKBUFX3 U5456 ( .A(n6380), .Y(n6373) );
  CLKBUFX3 U5457 ( .A(n6292), .Y(n6354) );
  CLKBUFX3 U5458 ( .A(n6292), .Y(n6356) );
  CLKBUFX3 U5459 ( .A(n6380), .Y(n6375) );
  CLKBUFX3 U5460 ( .A(n6292), .Y(n6355) );
  CLKBUFX3 U5461 ( .A(n6379), .Y(n6377) );
  CLKBUFX3 U5462 ( .A(n5744), .Y(n6304) );
  NAND2X1 U5463 ( .A(n6373), .B(n6472), .Y(n5744) );
  CLKINVX1 U5464 ( .A(n5632), .Y(n4574) );
  CLKINVX1 U5465 ( .A(n5840), .Y(n4593) );
  CLKINVX1 U5466 ( .A(n5644), .Y(n4588) );
  CLKINVX1 U5467 ( .A(n5610), .Y(n4599) );
  CLKINVX1 U5468 ( .A(n5642), .Y(n4598) );
  CLKINVX1 U5469 ( .A(n5608), .Y(n4589) );
  CLKINVX1 U5470 ( .A(n5645), .Y(n4568) );
  CLKINVX1 U5471 ( .A(n5611), .Y(n4569) );
  CLKINVX1 U5472 ( .A(n5612), .Y(n4563) );
  CLKINVX1 U5473 ( .A(n5183), .Y(n4573) );
  CLKINVX1 U5474 ( .A(n5246), .Y(n4584) );
  CLKINVX1 U5475 ( .A(n5248), .Y(n4562) );
  INVX3 U5476 ( .A(n6294), .Y(n6296) );
  INVX3 U5477 ( .A(n6294), .Y(n6297) );
  CLKINVX1 U5478 ( .A(n5082), .Y(n4508) );
  CLKINVX1 U5479 ( .A(n5126), .Y(n4553) );
  CLKBUFX3 U5480 ( .A(n6379), .Y(n6378) );
  NAND2X1 U5481 ( .A(n4511), .B(n4648), .Y(n5131) );
  CLKINVX1 U5482 ( .A(n5342), .Y(n4565) );
  CLKINVX1 U5483 ( .A(n5570), .Y(n4570) );
  CLKINVX1 U5484 ( .A(n5884), .Y(n4583) );
  CLKINVX1 U5485 ( .A(n5568), .Y(n4564) );
  CLKINVX1 U5486 ( .A(n5571), .Y(n4590) );
  CLKINVX1 U5487 ( .A(n5518), .Y(n4571) );
  CLKINVX1 U5488 ( .A(n5484), .Y(n4516) );
  CLKINVX1 U5489 ( .A(n5262), .Y(n4596) );
  CLKINVX1 U5490 ( .A(n5172), .Y(n4592) );
  CLKINVX1 U5491 ( .A(n5272), .Y(n4578) );
  CLKINVX1 U5492 ( .A(n5261), .Y(n4586) );
  NOR3X1 U5493 ( .A(n5150), .B(n5151), .C(n5152), .Y(n5142) );
  CLKINVX1 U5494 ( .A(n5257), .Y(n4600) );
  CLKBUFX3 U5495 ( .A(n5580), .Y(n6303) );
  INVX3 U5496 ( .A(n6294), .Y(n6295) );
  CLKINVX1 U5497 ( .A(n5337), .Y(n4575) );
  CLKINVX1 U5498 ( .A(n5127), .Y(n4556) );
  CLKBUFX3 U5499 ( .A(n5576), .Y(n6382) );
  CLKBUFX3 U5500 ( .A(n5574), .Y(n6384) );
  INVX3 U5501 ( .A(n5927), .Y(n4863) );
  CLKBUFX3 U5502 ( .A(n6380), .Y(n6376) );
  CLKINVX1 U5503 ( .A(n5441), .Y(n4551) );
  CLKINVX1 U5504 ( .A(n5444), .Y(n4546) );
  CLKBUFX3 U5505 ( .A(n6410), .Y(n6447) );
  CLKBUFX3 U5506 ( .A(n6410), .Y(n6446) );
  CLKBUFX3 U5507 ( .A(n6410), .Y(n6445) );
  CLKBUFX3 U5508 ( .A(n6411), .Y(n6450) );
  CLKBUFX3 U5509 ( .A(n6411), .Y(n6449) );
  CLKBUFX3 U5510 ( .A(n6411), .Y(n6448) );
  CLKBUFX3 U5511 ( .A(n6408), .Y(n6439) );
  CLKBUFX3 U5512 ( .A(n6409), .Y(n6444) );
  CLKBUFX3 U5513 ( .A(n6409), .Y(n6443) );
  CLKBUFX3 U5514 ( .A(n6409), .Y(n6442) );
  CLKBUFX3 U5515 ( .A(n6408), .Y(n6441) );
  CLKBUFX3 U5516 ( .A(n6408), .Y(n6440) );
  INVX3 U5517 ( .A(n6319), .Y(n4428) );
  INVX3 U5518 ( .A(n6318), .Y(n4427) );
  INVX3 U5519 ( .A(n6329), .Y(n4438) );
  INVX3 U5520 ( .A(n6328), .Y(n4437) );
  INVX3 U5521 ( .A(n6325), .Y(n4434) );
  INVX3 U5522 ( .A(n6324), .Y(n4433) );
  INVX3 U5523 ( .A(n6321), .Y(n4430) );
  INVX3 U5524 ( .A(n6320), .Y(n4429) );
  INVX3 U5525 ( .A(n6331), .Y(n4439) );
  INVX3 U5526 ( .A(n6327), .Y(n4436) );
  INVX3 U5527 ( .A(n6326), .Y(n4435) );
  INVX3 U5528 ( .A(n6323), .Y(n4432) );
  INVX3 U5529 ( .A(n6322), .Y(n4431) );
  INVX3 U5530 ( .A(n6341), .Y(n4446) );
  INVX3 U5531 ( .A(n6340), .Y(n4445) );
  INVX3 U5532 ( .A(n6337), .Y(n4442) );
  INVX3 U5533 ( .A(n6336), .Y(n4441) );
  INVX3 U5534 ( .A(n6342), .Y(n4447) );
  INVX3 U5535 ( .A(n6339), .Y(n4444) );
  INVX3 U5536 ( .A(n6338), .Y(n4443) );
  INVX3 U5537 ( .A(n6334), .Y(n4440) );
  INVX3 U5538 ( .A(n6347), .Y(n4448) );
  CLKBUFX3 U5539 ( .A(n5022), .Y(n6310) );
  OAI31XL U5540 ( .A0(n5037), .A1(n5035), .A2(n5036), .B0(n6308), .Y(n5022) );
  CLKBUFX3 U5541 ( .A(n5021), .Y(n6311) );
  OAI31XL U5542 ( .A0(n5037), .A1(n5036), .A2(n6290), .B0(n6308), .Y(n5021) );
  CLKBUFX3 U5543 ( .A(n5023), .Y(n6309) );
  OAI31XL U5544 ( .A0(n5037), .A1(n6290), .A2(n4544), .B0(n6308), .Y(n5023) );
  CLKBUFX3 U5545 ( .A(n5020), .Y(n6312) );
  OAI31XL U5546 ( .A0(n4544), .A1(n5035), .A2(n5034), .B0(n6308), .Y(n5020) );
  INVX16 U5547 ( .A(n6476), .Y(match_index[3]) );
  NAND4X1 U5548 ( .A(n5289), .B(n5290), .C(n5291), .D(n5292), .Y(n5086) );
  XNOR2X1 U5549 ( .A(n5251), .B(n5245), .Y(n5290) );
  XOR2X1 U5550 ( .A(n5244), .B(n4574), .Y(n5289) );
  NOR4X1 U5551 ( .A(n5293), .B(n5294), .C(n5295), .D(n5296), .Y(n5292) );
  XNOR2X1 U5552 ( .A(n5369), .B(n5363), .Y(n5402) );
  XNOR2X1 U5553 ( .A(n5374), .B(n5359), .Y(n5400) );
  XOR2X1 U5554 ( .A(n5373), .B(n5361), .Y(n5401) );
  XOR2X1 U5555 ( .A(n5384), .B(n5350), .Y(n5399) );
  NAND4X1 U5556 ( .A(n5313), .B(n5314), .C(n5315), .D(n5316), .Y(n5126) );
  XOR2X1 U5557 ( .A(n5335), .B(n4585), .Y(n5314) );
  XOR2X1 U5558 ( .A(n5336), .B(n4561), .Y(n5313) );
  NOR4X1 U5559 ( .A(n5317), .B(n5318), .C(n5319), .D(n5320), .Y(n5316) );
  NAND2X1 U5560 ( .A(n4457), .B(n4469), .Y(n4916) );
  NAND4X1 U5561 ( .A(n5395), .B(n5396), .C(n5397), .D(n5398), .Y(n5127) );
  XOR2X1 U5562 ( .A(n5352), .B(n4614), .Y(n5396) );
  XOR2X1 U5563 ( .A(n5354), .B(n4639), .Y(n5395) );
  NOR4X1 U5564 ( .A(n5399), .B(n5400), .C(n5401), .D(n5402), .Y(n5398) );
  NOR4X1 U5565 ( .A(n5412), .B(n5413), .C(n5414), .D(n5415), .Y(n5411) );
  XOR2X1 U5566 ( .A(n5360), .B(n5421), .Y(n5412) );
  XOR2X1 U5567 ( .A(n5364), .B(n5420), .Y(n5413) );
  XOR2X1 U5568 ( .A(n5351), .B(n5419), .Y(n5414) );
  NAND2X1 U5569 ( .A(n4912), .B(n6308), .Y(n4913) );
  XOR2X1 U5570 ( .A(n5331), .B(n5332), .Y(n5330) );
  CLKINVX1 U5571 ( .A(n6308), .Y(n4457) );
  XOR2X1 U5572 ( .A(n5232), .B(n4593), .Y(n5311) );
  XOR2X1 U5573 ( .A(n5337), .B(n4576), .Y(n5312) );
  NAND2X1 U5574 ( .A(n5067), .B(n5045), .Y(n5068) );
  CLKBUFX3 U5575 ( .A(n4969), .Y(n6316) );
  NAND2X1 U5576 ( .A(n4966), .B(n4931), .Y(n4969) );
  CLKBUFX3 U5577 ( .A(n4947), .Y(n6332) );
  NAND2X1 U5578 ( .A(n4944), .B(n4931), .Y(n4947) );
  XOR2X1 U5579 ( .A(n5350), .B(n5351), .Y(n5147) );
  XOR2X1 U5580 ( .A(n5354), .B(n5355), .Y(n5144) );
  XOR2X1 U5581 ( .A(n5359), .B(n5360), .Y(n5150) );
  XOR2X1 U5582 ( .A(n5363), .B(n5364), .Y(n5151) );
  INVX16 U5583 ( .A(n6454), .Y(match_index[0]) );
  XOR2X1 U5584 ( .A(n5352), .B(n5353), .Y(n5146) );
  XOR2X1 U5585 ( .A(n5361), .B(n5362), .Y(n5152) );
  NOR2X2 U5586 ( .A(n6463), .B(match_index[0]), .Y(n5701) );
  OAI22X1 U5587 ( .A0(n6455), .A1(n5681), .B0(n6296), .B1(n5682), .Y(n5327) );
  OAI22X1 U5588 ( .A0(n6456), .A1(n5813), .B0(n6296), .B1(n5778), .Y(n5240) );
  OAI22X1 U5589 ( .A0(n6455), .A1(n5658), .B0(n6295), .B1(n5674), .Y(n5331) );
  NOR4X1 U5590 ( .A(n5148), .B(n5144), .C(n5146), .D(n5147), .Y(n5349) );
  NOR4X1 U5591 ( .A(n5689), .B(n5690), .C(n5691), .D(n5692), .Y(n5688) );
  CLKINVX1 U5592 ( .A(n5383), .Y(n4614) );
  NAND4X1 U5593 ( .A(n5192), .B(n5193), .C(n5194), .D(n5195), .Y(n5134) );
  XNOR2X1 U5594 ( .A(n5251), .B(n5252), .Y(n5193) );
  XOR2X1 U5595 ( .A(n5253), .B(n4574), .Y(n5192) );
  NOR4X1 U5596 ( .A(n5196), .B(n5197), .C(n5198), .D(n5199), .Y(n5195) );
  CLKINVX1 U5597 ( .A(n5384), .Y(n4608) );
  CLKINVX1 U5598 ( .A(n5373), .Y(n4632) );
  NOR3X1 U5599 ( .A(n5174), .B(n4648), .C(n5138), .Y(n5159) );
  XOR2X1 U5600 ( .A(n4578), .B(n4505), .Y(n5174) );
  NOR3X1 U5601 ( .A(n5222), .B(n5223), .C(n5136), .Y(n5211) );
  XOR2X1 U5602 ( .A(n5245), .B(n4593), .Y(n5222) );
  XOR2X1 U5603 ( .A(n5244), .B(n4575), .Y(n5223) );
  CLKINVX1 U5604 ( .A(n5129), .Y(n4510) );
  OAI32X1 U5605 ( .A0(n5130), .A1(n5131), .A2(n5085), .B0(n4648), .B1(n5132), 
        .Y(n5129) );
  CLKBUFX3 U5606 ( .A(n6468), .Y(n6473) );
  CLKBUFX3 U5607 ( .A(n5702), .Y(n6357) );
  OAI32X1 U5608 ( .A0(n5135), .A1(n5126), .A2(n5131), .B0(n4648), .B1(n5136), 
        .Y(n5082) );
  OAI22X1 U5609 ( .A0(n6455), .A1(n5622), .B0(n6296), .B1(n5653), .Y(n5248) );
  NAND2X2 U5610 ( .A(n4554), .B(n5372), .Y(n5370) );
  OAI22X1 U5611 ( .A0(n6456), .A1(n5542), .B0(n6295), .B1(n5635), .Y(n5183) );
  OAI22X1 U5612 ( .A0(n6456), .A1(n5849), .B0(n6296), .B1(n5813), .Y(n5246) );
  AOI222XL U5613 ( .A0(n4542), .A1(n4556), .B0(n4547), .B1(n4609), .C0(n4548), 
        .C1(n4553), .Y(n5074) );
  XNOR2X1 U5614 ( .A(n5375), .B(n5322), .Y(n5365) );
  XOR2X1 U5615 ( .A(n5382), .B(n5332), .Y(n5379) );
  XOR2X1 U5616 ( .A(n5383), .B(n5324), .Y(n5378) );
  XOR2X1 U5617 ( .A(n5384), .B(n5334), .Y(n5377) );
  OA22X1 U5618 ( .A0(n6458), .A1(n5870), .B0(n6295), .B1(n5849), .Y(n5204) );
  OA22X1 U5619 ( .A0(n6458), .A1(n5857), .B0(n6296), .B1(n5681), .Y(n5221) );
  OA22X1 U5620 ( .A0(n6458), .A1(n5599), .B0(n6296), .B1(n5857), .Y(n5202) );
  XOR2X1 U5621 ( .A(n5183), .B(n5253), .Y(n5284) );
  XOR2X1 U5622 ( .A(n5373), .B(n5336), .Y(n5367) );
  OA22X1 U5623 ( .A0(n6458), .A1(n5864), .B0(n6295), .B1(n5843), .Y(n5251) );
  XOR2X1 U5624 ( .A(n5220), .B(n5202), .Y(n5295) );
  XOR2X1 U5625 ( .A(n5247), .B(n5204), .Y(n5294) );
  XOR2X1 U5626 ( .A(n5234), .B(n5221), .Y(n5305) );
  NAND2X2 U5627 ( .A(n4554), .B(n5149), .Y(n5372) );
  XOR2X1 U5628 ( .A(n5232), .B(n4594), .Y(n5231) );
  XOR2X1 U5629 ( .A(n5234), .B(n4581), .Y(n5228) );
  XOR2X1 U5630 ( .A(n4577), .B(n4576), .Y(n5229) );
  AO22X1 U5631 ( .A0(n5636), .A1(n6296), .B0(n6457), .B1(n5819), .Y(n5337) );
  CLKINVX1 U5632 ( .A(n5344), .Y(n4507) );
  CLKBUFX3 U5633 ( .A(n6468), .Y(n6474) );
  CLKINVX1 U5634 ( .A(n5085), .Y(n4552) );
  CLKINVX1 U5635 ( .A(n6454), .Y(n6453) );
  CLKBUFX3 U5636 ( .A(n6459), .Y(n6457) );
  OAI22X1 U5637 ( .A0(n6456), .A1(n5531), .B0(n6295), .B1(n5590), .Y(n5257) );
  NAND4X1 U5638 ( .A(n5133), .B(n5137), .C(n5155), .D(n5489), .Y(n5484) );
  AND3X2 U5639 ( .A(n5135), .B(n5130), .C(n5345), .Y(n5489) );
  XNOR2X1 U5640 ( .A(match_index[1]), .B(n5452), .Y(n5386) );
  OAI22X1 U5641 ( .A0(n6454), .A1(n5510), .B0(n6297), .B1(n5542), .Y(n5272) );
  OAI22X1 U5642 ( .A0(n6454), .A1(n5521), .B0(match_index[0]), .B1(n5522), .Y(
        n5261) );
  OAI22X1 U5643 ( .A0(match_index[0]), .A1(n5548), .B0(n6456), .B1(n5549), .Y(
        n5172) );
  XOR2X1 U5644 ( .A(n5272), .B(n5184), .Y(n5271) );
  XOR2X1 U5645 ( .A(n5183), .B(n5184), .Y(n5182) );
  OA22X1 U5646 ( .A0(n6458), .A1(n5548), .B0(n6295), .B1(n5864), .Y(n5187) );
  OA22X1 U5647 ( .A0(n6458), .A1(n5554), .B0(n6295), .B1(n5555), .Y(n5165) );
  OA22X1 U5648 ( .A0(n6458), .A1(n5539), .B0(n6297), .B1(n5540), .Y(n5173) );
  OA22X1 U5649 ( .A0(n6458), .A1(n5555), .B0(n6297), .B1(n5599), .Y(n5255) );
  XOR2X1 U5650 ( .A(n5201), .B(n5202), .Y(n5198) );
  XOR2X1 U5651 ( .A(n5252), .B(n5187), .Y(n5282) );
  XOR2X1 U5652 ( .A(n5203), .B(n5204), .Y(n5197) );
  XOR2X1 U5653 ( .A(n5186), .B(n5187), .Y(n5180) );
  XOR2X1 U5654 ( .A(n5220), .B(n5221), .Y(n5213) );
  XOR2X1 U5655 ( .A(n5186), .B(n4592), .Y(n5268) );
  XOR2X1 U5656 ( .A(n4579), .B(n4505), .Y(n5106) );
  NOR4X1 U5657 ( .A(n5144), .B(n5145), .C(n5146), .D(n5147), .Y(n5143) );
  NAND2BX1 U5658 ( .AN(n5148), .B(n5149), .Y(n5145) );
  XNOR2X1 U5659 ( .A(n5173), .B(n5124), .Y(n5170) );
  CLKINVX1 U5660 ( .A(n5472), .Y(n4515) );
  CLKINVX1 U5661 ( .A(n5067), .Y(n4511) );
  CLKBUFX3 U5662 ( .A(n6458), .Y(n6455) );
  CLKBUFX3 U5663 ( .A(n6458), .Y(n6456) );
  CLKBUFX3 U5664 ( .A(n6459), .Y(n6458) );
  XOR2X1 U5665 ( .A(n5393), .B(n5456), .Y(n5450) );
  XOR2X1 U5666 ( .A(n6473), .B(n5452), .Y(n5456) );
  XOR2X1 U5667 ( .A(match_index[3]), .B(n5453), .Y(n5451) );
  NAND2X1 U5668 ( .A(n5454), .B(n5455), .Y(n5453) );
  OAI21XL U5669 ( .A0(n5393), .A1(n5452), .B0(n4513), .Y(n5455) );
  XOR2X1 U5670 ( .A(n5172), .B(n5117), .Y(n5171) );
  NAND2X1 U5671 ( .A(n4648), .B(n5067), .Y(n5075) );
  OR3X2 U5672 ( .A(n5452), .B(n4513), .C(n5393), .Y(n5454) );
  NAND2X1 U5673 ( .A(n4506), .B(n5454), .Y(n5470) );
  OAI21XL U5674 ( .A0(n4506), .A1(n5454), .B0(n5470), .Y(n5480) );
  INVX3 U5675 ( .A(n5149), .Y(n4648) );
  XOR2X1 U5676 ( .A(n5040), .B(n4550), .Y(n5436) );
  XOR2X1 U5677 ( .A(n5091), .B(n5924), .Y(n5441) );
  NAND2X1 U5678 ( .A(n4551), .B(n5056), .Y(n5444) );
  CLKINVX1 U5679 ( .A(n4987), .Y(n4829) );
  CLKINVX1 U5680 ( .A(n5926), .Y(n4550) );
  CLKINVX1 U5681 ( .A(n5080), .Y(n4547) );
  CLKINVX1 U5682 ( .A(n5056), .Y(n4545) );
  CLKINVX1 U5683 ( .A(n4992), .Y(n4830) );
  XNOR2X1 U5684 ( .A(n5091), .B(n5088), .Y(n5039) );
  CLKBUFX3 U5685 ( .A(n6412), .Y(n6410) );
  CLKBUFX3 U5686 ( .A(n6444), .Y(n6411) );
  CLKBUFX3 U5687 ( .A(n6413), .Y(n6407) );
  CLKBUFX3 U5688 ( .A(n6412), .Y(n6409) );
  CLKBUFX3 U5689 ( .A(n6413), .Y(n6408) );
  OAI22XL U5690 ( .A0(n6033), .A1(n5026), .B0(n4456), .B1(n5027), .Y(n1366) );
  OAI22XL U5691 ( .A0(n6032), .A1(n5026), .B0(n4456), .B1(n5028), .Y(n1359) );
  OAI22XL U5692 ( .A0(n6034), .A1(n5026), .B0(n4456), .B1(n5029), .Y(n1352) );
  OAI22XL U5693 ( .A0(n6013), .A1(n5026), .B0(n4456), .B1(n5030), .Y(n1345) );
  OAI22XL U5694 ( .A0(n6014), .A1(n5026), .B0(n4456), .B1(n5031), .Y(n1338) );
  OAI22XL U5695 ( .A0(n5985), .A1(n5026), .B0(n4456), .B1(n5032), .Y(n1331) );
  OAI22XL U5696 ( .A0(n6298), .A1(n4978), .B0(n4999), .B1(n6020), .Y(n1397) );
  OAI22XL U5697 ( .A0(n6298), .A1(n4984), .B0(n6056), .B1(n4999), .Y(n1392) );
  OAI22XL U5698 ( .A0(n6298), .A1(n4981), .B0(n6065), .B1(n4999), .Y(n1395) );
  OAI22XL U5699 ( .A0(n6298), .A1(n4982), .B0(n5987), .B1(n4999), .Y(n1394) );
  OAI22XL U5700 ( .A0(n6298), .A1(n4979), .B0(n6025), .B1(n4999), .Y(n1396) );
  NAND3X1 U5701 ( .A(n5038), .B(n5039), .C(n6006), .Y(n5034) );
  OAI21X2 U5702 ( .A0(n4987), .A1(n4988), .B0(n4989), .Y(n4980) );
  OAI21X2 U5703 ( .A0(n4974), .A1(n4997), .B0(n4989), .Y(n5000) );
  OAI21X2 U5704 ( .A0(n4995), .A1(n4993), .B0(n4989), .Y(n4994) );
  OAI21X2 U5705 ( .A0(n4987), .A1(n4997), .B0(n4989), .Y(n4996) );
  OAI21X2 U5706 ( .A0(n4973), .A1(n4997), .B0(n4989), .Y(n4998) );
  NOR2BX1 U5707 ( .AN(n4948), .B(n4851), .Y(n4954) );
  CLKBUFX3 U5708 ( .A(n4914), .Y(n6313) );
  NAND3BX1 U5709 ( .AN(next_state[1]), .B(next_state[0]), .C(n5014), .Y(n4914)
         );
  OAI22XL U5710 ( .A0(n5981), .A1(n5019), .B0(n6300), .B1(n5018), .Y(n1372) );
  OAI22XL U5711 ( .A0(n5996), .A1(n5019), .B0(n6300), .B1(n5030), .Y(n1343) );
  OAI22XL U5712 ( .A0(n5979), .A1(n5019), .B0(n6300), .B1(n5032), .Y(n1329) );
  OAI22XL U5713 ( .A0(n6300), .A1(n5033), .B0(n6037), .B1(n5019), .Y(n1322) );
  CLKBUFX3 U5714 ( .A(n4990), .Y(n6315) );
  OAI21XL U5715 ( .A0(n4973), .A1(n4988), .B0(n4989), .Y(n4990) );
  CLKBUFX3 U5716 ( .A(n4991), .Y(n6314) );
  OAI21XL U5717 ( .A0(n4992), .A1(n4993), .B0(n4989), .Y(n4991) );
  OAI22XL U5718 ( .A0(n5000), .A1(n6017), .B0(n4459), .B1(n4978), .Y(n1389) );
  OAI22XL U5719 ( .A0(n6063), .A1(n5000), .B0(n4459), .B1(n4984), .Y(n1384) );
  OAI22XL U5720 ( .A0(n6070), .A1(n5000), .B0(n4459), .B1(n4981), .Y(n1387) );
  OAI22XL U5721 ( .A0(n5989), .A1(n5000), .B0(n4459), .B1(n4982), .Y(n1386) );
  OAI22XL U5722 ( .A0(n6026), .A1(n5000), .B0(n4459), .B1(n4979), .Y(n1388) );
  OAI22XL U5723 ( .A0(n4464), .A1(n4979), .B0(n6015), .B1(n4980), .Y(n1444) );
  OAI22XL U5724 ( .A0(n4464), .A1(n4981), .B0(n6031), .B1(n4980), .Y(n1443) );
  OAI22XL U5725 ( .A0(n4464), .A1(n4982), .B0(n6016), .B1(n4980), .Y(n1442) );
  OAI22XL U5726 ( .A0(n4464), .A1(n4983), .B0(n6010), .B1(n4980), .Y(n1441) );
  OAI22XL U5727 ( .A0(n4464), .A1(n4984), .B0(n6008), .B1(n4980), .Y(n1440) );
  OAI22XL U5728 ( .A0(n4464), .A1(n4985), .B0(n5983), .B1(n4980), .Y(n1439) );
  OAI22XL U5729 ( .A0(n4466), .A1(n4978), .B0(n4994), .B1(n4871), .Y(n1421) );
  OAI22XL U5730 ( .A0(n4462), .A1(n4978), .B0(n4996), .B1(n6018), .Y(n1413) );
  OAI22XL U5731 ( .A0(n4461), .A1(n4978), .B0(n4998), .B1(n6019), .Y(n1405) );
  OAI22XL U5732 ( .A0(n6043), .A1(n6310), .B0(n4451), .B1(n5029), .Y(n1347) );
  OAI22XL U5733 ( .A0(n6044), .A1(n6310), .B0(n4451), .B1(n5030), .Y(n1340) );
  OAI22XL U5734 ( .A0(n6057), .A1(n6310), .B0(n4451), .B1(n5031), .Y(n1333) );
  OAI22XL U5735 ( .A0(n6055), .A1(n6310), .B0(n4451), .B1(n5032), .Y(n1326) );
  OAI22XL U5736 ( .A0(n5992), .A1(n6312), .B0(n4453), .B1(n5027), .Y(n1363) );
  OAI22XL U5737 ( .A0(n6042), .A1(n6312), .B0(n4453), .B1(n5028), .Y(n1357) );
  OAI22XL U5738 ( .A0(n6035), .A1(n6312), .B0(n4453), .B1(n5029), .Y(n1349) );
  OAI22XL U5739 ( .A0(n5997), .A1(n6312), .B0(n4453), .B1(n5030), .Y(n1342) );
  OAI22XL U5740 ( .A0(n6041), .A1(n6312), .B0(n4453), .B1(n5031), .Y(n1335) );
  OAI22XL U5741 ( .A0(n6039), .A1(n6312), .B0(n4453), .B1(n5032), .Y(n1328) );
  OAI22XL U5742 ( .A0(n5990), .A1(n6312), .B0(n4453), .B1(n5018), .Y(n1371) );
  OAI22XL U5743 ( .A0(n5993), .A1(n6311), .B0(n4452), .B1(n5018), .Y(n1370) );
  OAI22XL U5744 ( .A0(n5995), .A1(n6310), .B0(n4451), .B1(n5018), .Y(n1369) );
  OAI22XL U5745 ( .A0(n6036), .A1(n6311), .B0(n4452), .B1(n5029), .Y(n1348) );
  OAI22XL U5746 ( .A0(n5994), .A1(n6311), .B0(n4452), .B1(n5027), .Y(n1362) );
  OAI22XL U5747 ( .A0(n5998), .A1(n6310), .B0(n4451), .B1(n5027), .Y(n1361) );
  OAI22XL U5748 ( .A0(n6038), .A1(n6311), .B0(n4452), .B1(n5030), .Y(n1341) );
  OAI22XL U5749 ( .A0(n6045), .A1(n6311), .B0(n4452), .B1(n5032), .Y(n1327) );
  OAI22XL U5750 ( .A0(n6049), .A1(n6311), .B0(n4452), .B1(n5031), .Y(n1334) );
  OAI22XL U5751 ( .A0(n6050), .A1(n6311), .B0(n4452), .B1(n5028), .Y(n1356) );
  OAI22XL U5752 ( .A0(n6058), .A1(n6310), .B0(n4451), .B1(n5028), .Y(n1355) );
  OAI22XL U5753 ( .A0(n6061), .A1(n6309), .B0(n4450), .B1(n5030), .Y(n1339) );
  OAI22XL U5754 ( .A0(n6002), .A1(n6309), .B0(n4450), .B1(n5032), .Y(n1325) );
  OAI22XL U5755 ( .A0(n6054), .A1(n6309), .B0(n4450), .B1(n5033), .Y(n1318) );
  OAI22XL U5756 ( .A0(n5999), .A1(n6309), .B0(n4450), .B1(n5018), .Y(n1368) );
  OAI22XL U5757 ( .A0(n6053), .A1(n6309), .B0(n4450), .B1(n5029), .Y(n1346) );
  OAI22XL U5758 ( .A0(n6001), .A1(n6309), .B0(n4450), .B1(n5027), .Y(n1360) );
  OAI22XL U5759 ( .A0(n6062), .A1(n6309), .B0(n4450), .B1(n5031), .Y(n1332) );
  OAI22XL U5760 ( .A0(n6064), .A1(n6309), .B0(n4450), .B1(n5028), .Y(n1354) );
  OAI22XL U5761 ( .A0(n4466), .A1(n4979), .B0(n4870), .B1(n4994), .Y(n1420) );
  OAI22XL U5762 ( .A0(n4466), .A1(n4981), .B0(n4869), .B1(n4994), .Y(n1419) );
  OAI22XL U5763 ( .A0(n4466), .A1(n4982), .B0(n4868), .B1(n4994), .Y(n1418) );
  OAI22XL U5764 ( .A0(n4466), .A1(n4984), .B0(n4867), .B1(n4994), .Y(n1416) );
  OAI22XL U5765 ( .A0(n4462), .A1(n4982), .B0(n5986), .B1(n4996), .Y(n1410) );
  OAI22XL U5766 ( .A0(n4462), .A1(n4979), .B0(n6023), .B1(n4996), .Y(n1412) );
  OAI22XL U5767 ( .A0(n4462), .A1(n4984), .B0(n6047), .B1(n4996), .Y(n1408) );
  OAI22XL U5768 ( .A0(n4461), .A1(n4984), .B0(n6048), .B1(n4998), .Y(n1400) );
  OAI22XL U5769 ( .A0(n4462), .A1(n4981), .B0(n6051), .B1(n4996), .Y(n1411) );
  OAI22XL U5770 ( .A0(n4461), .A1(n4981), .B0(n6059), .B1(n4998), .Y(n1403) );
  OAI22XL U5771 ( .A0(n4461), .A1(n4982), .B0(n5988), .B1(n4998), .Y(n1402) );
  OAI22XL U5772 ( .A0(n4461), .A1(n4979), .B0(n6024), .B1(n4998), .Y(n1404) );
  OAI22XL U5773 ( .A0(n4463), .A1(n4986), .B0(n6315), .B1(n6029), .Y(n1430) );
  OAI22XL U5774 ( .A0(n4467), .A1(n4986), .B0(n6314), .B1(n4872), .Y(n1422) );
  OAI22XL U5775 ( .A0(n4463), .A1(n4983), .B0(n6315), .B1(n6030), .Y(n1433) );
  OAI22XL U5776 ( .A0(n4463), .A1(n4985), .B0(n6315), .B1(n6028), .Y(n1431) );
  OAI22XL U5777 ( .A0(n4467), .A1(n4983), .B0(n6314), .B1(n4874), .Y(n1425) );
  OAI22XL U5778 ( .A0(n4467), .A1(n4985), .B0(n6314), .B1(n4873), .Y(n1423) );
  OAI22XL U5779 ( .A0(n4463), .A1(n4978), .B0(n6315), .B1(n6027), .Y(n1437) );
  OAI22XL U5780 ( .A0(n4467), .A1(n4979), .B0(n4878), .B1(n6314), .Y(n1428) );
  OAI22XL U5781 ( .A0(n4467), .A1(n4981), .B0(n4877), .B1(n6314), .Y(n1427) );
  OAI22XL U5782 ( .A0(n4467), .A1(n4982), .B0(n4876), .B1(n6314), .Y(n1426) );
  OAI22XL U5783 ( .A0(n4467), .A1(n4984), .B0(n4875), .B1(n6314), .Y(n1424) );
  OAI22XL U5784 ( .A0(n4428), .A1(n4827), .B0(n6391), .B1(n6319), .Y(n1483) );
  OAI22XL U5785 ( .A0(n4428), .A1(n4826), .B0(n6394), .B1(n6319), .Y(n1482) );
  OAI22XL U5786 ( .A0(n4428), .A1(n4825), .B0(n6395), .B1(n6319), .Y(n1481) );
  OAI22XL U5787 ( .A0(n4428), .A1(n4824), .B0(n6397), .B1(n6319), .Y(n1480) );
  OAI22XL U5788 ( .A0(n4428), .A1(n4823), .B0(n6399), .B1(n6319), .Y(n1479) );
  OAI22XL U5789 ( .A0(n4428), .A1(n4822), .B0(n6401), .B1(n6319), .Y(n1478) );
  OAI22XL U5790 ( .A0(n4428), .A1(n4821), .B0(n6403), .B1(n6319), .Y(n1477) );
  OAI22XL U5791 ( .A0(n4428), .A1(n4820), .B0(n6405), .B1(n6319), .Y(n1476) );
  OAI22XL U5792 ( .A0(n4427), .A1(n4819), .B0(n6391), .B1(n6318), .Y(n1475) );
  OAI22XL U5793 ( .A0(n4427), .A1(n4818), .B0(n6393), .B1(n6318), .Y(n1474) );
  OAI22XL U5794 ( .A0(n4427), .A1(n4817), .B0(n6395), .B1(n6318), .Y(n1473) );
  OAI22XL U5795 ( .A0(n4427), .A1(n4816), .B0(n6397), .B1(n6318), .Y(n1472) );
  OAI22XL U5796 ( .A0(n4427), .A1(n4815), .B0(n6399), .B1(n6318), .Y(n1471) );
  OAI22XL U5797 ( .A0(n4427), .A1(n4814), .B0(n6401), .B1(n6318), .Y(n1470) );
  OAI22XL U5798 ( .A0(n4427), .A1(n4813), .B0(n6403), .B1(n6318), .Y(n1469) );
  OAI22XL U5799 ( .A0(n4427), .A1(n4812), .B0(n6405), .B1(n6318), .Y(n1468) );
  OAI22XL U5800 ( .A0(n4438), .A1(n4811), .B0(n6392), .B1(n6329), .Y(n1563) );
  OAI22XL U5801 ( .A0(n4438), .A1(n4810), .B0(n6394), .B1(n6329), .Y(n1562) );
  OAI22XL U5802 ( .A0(n4438), .A1(n4809), .B0(n6396), .B1(n6329), .Y(n1561) );
  OAI22XL U5803 ( .A0(n4438), .A1(n4808), .B0(n6398), .B1(n6329), .Y(n1560) );
  OAI22XL U5804 ( .A0(n4438), .A1(n4807), .B0(n6400), .B1(n6329), .Y(n1559) );
  OAI22XL U5805 ( .A0(n4438), .A1(n4806), .B0(n6402), .B1(n6329), .Y(n1558) );
  OAI22XL U5806 ( .A0(n4438), .A1(n4805), .B0(n6404), .B1(n6329), .Y(n1557) );
  OAI22XL U5807 ( .A0(n4438), .A1(n4804), .B0(n6406), .B1(n6329), .Y(n1556) );
  OAI22XL U5808 ( .A0(n4437), .A1(n4803), .B0(n6392), .B1(n6328), .Y(n1555) );
  OAI22XL U5809 ( .A0(n4437), .A1(n4802), .B0(n6394), .B1(n6328), .Y(n1554) );
  OAI22XL U5810 ( .A0(n4437), .A1(n4801), .B0(n6396), .B1(n6328), .Y(n1553) );
  OAI22XL U5811 ( .A0(n4437), .A1(n4800), .B0(n6398), .B1(n6328), .Y(n1552) );
  OAI22XL U5812 ( .A0(n4437), .A1(n4799), .B0(n6400), .B1(n6328), .Y(n1551) );
  OAI22XL U5813 ( .A0(n4437), .A1(n4798), .B0(n6402), .B1(n6328), .Y(n1550) );
  OAI22XL U5814 ( .A0(n4437), .A1(n4797), .B0(n6404), .B1(n6328), .Y(n1549) );
  OAI22XL U5815 ( .A0(n4437), .A1(n4796), .B0(n6406), .B1(n6328), .Y(n1548) );
  OAI22XL U5816 ( .A0(n4434), .A1(n4795), .B0(n6392), .B1(n6325), .Y(n1531) );
  OAI22XL U5817 ( .A0(n4434), .A1(n4794), .B0(n6394), .B1(n6325), .Y(n1530) );
  OAI22XL U5818 ( .A0(n4434), .A1(n4793), .B0(n6396), .B1(n6325), .Y(n1529) );
  OAI22XL U5819 ( .A0(n4434), .A1(n4792), .B0(n6398), .B1(n6325), .Y(n1528) );
  OAI22XL U5820 ( .A0(n4434), .A1(n4791), .B0(n6400), .B1(n6325), .Y(n1527) );
  OAI22XL U5821 ( .A0(n4434), .A1(n4790), .B0(n6402), .B1(n6325), .Y(n1526) );
  OAI22XL U5822 ( .A0(n4434), .A1(n4789), .B0(n6404), .B1(n6325), .Y(n1525) );
  OAI22XL U5823 ( .A0(n4434), .A1(n4788), .B0(n6406), .B1(n6325), .Y(n1524) );
  OAI22XL U5824 ( .A0(n4433), .A1(n4787), .B0(n6392), .B1(n6324), .Y(n1523) );
  OAI22XL U5825 ( .A0(n4433), .A1(n4786), .B0(n6394), .B1(n6324), .Y(n1522) );
  OAI22XL U5826 ( .A0(n4433), .A1(n4785), .B0(n6396), .B1(n6324), .Y(n1521) );
  OAI22XL U5827 ( .A0(n4433), .A1(n4784), .B0(n6398), .B1(n6324), .Y(n1520) );
  OAI22XL U5828 ( .A0(n4433), .A1(n4783), .B0(n6400), .B1(n6324), .Y(n1519) );
  OAI22XL U5829 ( .A0(n4433), .A1(n4782), .B0(n6402), .B1(n6324), .Y(n1518) );
  OAI22XL U5830 ( .A0(n4433), .A1(n4781), .B0(n6404), .B1(n6324), .Y(n1517) );
  OAI22XL U5831 ( .A0(n4433), .A1(n4780), .B0(n6406), .B1(n6324), .Y(n1516) );
  OAI22XL U5832 ( .A0(n4430), .A1(n4779), .B0(n6391), .B1(n6321), .Y(n1499) );
  OAI22XL U5833 ( .A0(n4430), .A1(n4778), .B0(n6394), .B1(n6321), .Y(n1498) );
  OAI22XL U5834 ( .A0(n4430), .A1(n4777), .B0(n6395), .B1(n6321), .Y(n1497) );
  OAI22XL U5835 ( .A0(n4430), .A1(n4776), .B0(n6397), .B1(n6321), .Y(n1496) );
  OAI22XL U5836 ( .A0(n4430), .A1(n4775), .B0(n6399), .B1(n6321), .Y(n1495) );
  OAI22XL U5837 ( .A0(n4430), .A1(n4774), .B0(n6401), .B1(n6321), .Y(n1494) );
  OAI22XL U5838 ( .A0(n4430), .A1(n4773), .B0(n6403), .B1(n6321), .Y(n1493) );
  OAI22XL U5839 ( .A0(n4430), .A1(n4772), .B0(n6405), .B1(n6321), .Y(n1492) );
  OAI22XL U5840 ( .A0(n4429), .A1(n4771), .B0(n6392), .B1(n6320), .Y(n1491) );
  OAI22XL U5841 ( .A0(n4429), .A1(n4770), .B0(n6394), .B1(n6320), .Y(n1490) );
  OAI22XL U5842 ( .A0(n4429), .A1(n4769), .B0(n6396), .B1(n6320), .Y(n1489) );
  OAI22XL U5843 ( .A0(n4429), .A1(n4768), .B0(n6398), .B1(n6320), .Y(n1488) );
  OAI22XL U5844 ( .A0(n4429), .A1(n4767), .B0(n6400), .B1(n6320), .Y(n1487) );
  OAI22XL U5845 ( .A0(n4429), .A1(n4766), .B0(n6402), .B1(n6320), .Y(n1486) );
  OAI22XL U5846 ( .A0(n4429), .A1(n4765), .B0(n6404), .B1(n6320), .Y(n1485) );
  OAI22XL U5847 ( .A0(n4429), .A1(n4764), .B0(n6406), .B1(n6320), .Y(n1484) );
  OAI22XL U5848 ( .A0(n4439), .A1(n4763), .B0(n6392), .B1(n6331), .Y(n1579) );
  OAI22XL U5849 ( .A0(n4439), .A1(n6012), .B0(n6394), .B1(n6331), .Y(n1578) );
  OAI22XL U5850 ( .A0(n4439), .A1(n4761), .B0(n6396), .B1(n6331), .Y(n1577) );
  OAI22XL U5851 ( .A0(n4439), .A1(n4760), .B0(n6398), .B1(n6331), .Y(n1576) );
  OAI22XL U5852 ( .A0(n4439), .A1(n4759), .B0(n6400), .B1(n6331), .Y(n1575) );
  OAI22XL U5853 ( .A0(n4439), .A1(n4758), .B0(n6402), .B1(n6331), .Y(n1574) );
  OAI22XL U5854 ( .A0(n4439), .A1(n4757), .B0(n6404), .B1(n6331), .Y(n1573) );
  OAI22XL U5855 ( .A0(n4439), .A1(n4756), .B0(n6406), .B1(n6331), .Y(n1572) );
  OAI22XL U5856 ( .A0(n4436), .A1(n4755), .B0(n6392), .B1(n6327), .Y(n1547) );
  OAI22XL U5857 ( .A0(n4436), .A1(n4754), .B0(n6394), .B1(n6327), .Y(n1546) );
  OAI22XL U5858 ( .A0(n4436), .A1(n4753), .B0(n6396), .B1(n6327), .Y(n1545) );
  OAI22XL U5859 ( .A0(n4436), .A1(n4752), .B0(n6398), .B1(n6327), .Y(n1544) );
  OAI22XL U5860 ( .A0(n4436), .A1(n4751), .B0(n6400), .B1(n6327), .Y(n1543) );
  OAI22XL U5861 ( .A0(n4436), .A1(n4750), .B0(n6402), .B1(n6327), .Y(n1542) );
  OAI22XL U5862 ( .A0(n4436), .A1(n4749), .B0(n6404), .B1(n6327), .Y(n1541) );
  OAI22XL U5863 ( .A0(n4436), .A1(n4748), .B0(n6406), .B1(n6327), .Y(n1540) );
  OAI22XL U5864 ( .A0(n4435), .A1(n4747), .B0(n6392), .B1(n6326), .Y(n1539) );
  OAI22XL U5865 ( .A0(n4435), .A1(n4746), .B0(n6394), .B1(n6326), .Y(n1538) );
  OAI22XL U5866 ( .A0(n4435), .A1(n4745), .B0(n6396), .B1(n6326), .Y(n1537) );
  OAI22XL U5867 ( .A0(n4435), .A1(n4744), .B0(n6398), .B1(n6326), .Y(n1536) );
  OAI22XL U5868 ( .A0(n4435), .A1(n4743), .B0(n6400), .B1(n6326), .Y(n1535) );
  OAI22XL U5869 ( .A0(n4435), .A1(n4742), .B0(n6402), .B1(n6326), .Y(n1534) );
  OAI22XL U5870 ( .A0(n4435), .A1(n4741), .B0(n6404), .B1(n6326), .Y(n1533) );
  OAI22XL U5871 ( .A0(n4435), .A1(n4740), .B0(n6406), .B1(n6326), .Y(n1532) );
  OAI22XL U5872 ( .A0(n4432), .A1(n4739), .B0(n6392), .B1(n6323), .Y(n1515) );
  OAI22XL U5873 ( .A0(n4432), .A1(n4738), .B0(n6394), .B1(n6323), .Y(n1514) );
  OAI22XL U5874 ( .A0(n4432), .A1(n4737), .B0(n6396), .B1(n6323), .Y(n1513) );
  OAI22XL U5875 ( .A0(n4432), .A1(n4736), .B0(n4841), .B1(n6323), .Y(n1512) );
  OAI22XL U5876 ( .A0(n4432), .A1(n4735), .B0(n6400), .B1(n6323), .Y(n1511) );
  OAI22XL U5877 ( .A0(n4432), .A1(n4734), .B0(n4839), .B1(n6323), .Y(n1510) );
  OAI22XL U5878 ( .A0(n4432), .A1(n4733), .B0(n6404), .B1(n6323), .Y(n1509) );
  OAI22XL U5879 ( .A0(n4432), .A1(n4732), .B0(n6406), .B1(n6323), .Y(n1508) );
  OAI22XL U5880 ( .A0(n4431), .A1(n4731), .B0(n4844), .B1(n6322), .Y(n1507) );
  OAI22XL U5881 ( .A0(n4431), .A1(n4730), .B0(n6394), .B1(n6322), .Y(n1506) );
  OAI22XL U5882 ( .A0(n4431), .A1(n4729), .B0(n4842), .B1(n6322), .Y(n1505) );
  OAI22XL U5883 ( .A0(n4431), .A1(n4728), .B0(n4841), .B1(n6322), .Y(n1504) );
  OAI22XL U5884 ( .A0(n4431), .A1(n4727), .B0(n4840), .B1(n6322), .Y(n1503) );
  OAI22XL U5885 ( .A0(n4431), .A1(n4726), .B0(n6402), .B1(n6322), .Y(n1502) );
  OAI22XL U5886 ( .A0(n4431), .A1(n4725), .B0(n4838), .B1(n6322), .Y(n1501) );
  OAI22XL U5887 ( .A0(n4431), .A1(n4724), .B0(n4837), .B1(n6322), .Y(n1500) );
  OAI22XL U5888 ( .A0(n4446), .A1(n4723), .B0(n6392), .B1(n6341), .Y(n1659) );
  OAI22XL U5889 ( .A0(n4446), .A1(n6009), .B0(n6394), .B1(n6341), .Y(n1658) );
  OAI22XL U5890 ( .A0(n4446), .A1(n4721), .B0(n6396), .B1(n6341), .Y(n1657) );
  OAI22XL U5891 ( .A0(n4446), .A1(n4720), .B0(n6398), .B1(n6341), .Y(n1656) );
  OAI22XL U5892 ( .A0(n4446), .A1(n4719), .B0(n6400), .B1(n6341), .Y(n1655) );
  OAI22XL U5893 ( .A0(n4446), .A1(n4718), .B0(n6402), .B1(n6341), .Y(n1654) );
  OAI22XL U5894 ( .A0(n4446), .A1(n4717), .B0(n6404), .B1(n6341), .Y(n1653) );
  OAI22XL U5895 ( .A0(n4446), .A1(n4716), .B0(n6406), .B1(n6341), .Y(n1652) );
  OAI22XL U5896 ( .A0(n4445), .A1(n4715), .B0(n6391), .B1(n6340), .Y(n1651) );
  OAI22XL U5897 ( .A0(n4445), .A1(n5982), .B0(n6394), .B1(n6340), .Y(n1650) );
  OAI22XL U5898 ( .A0(n4445), .A1(n4713), .B0(n6395), .B1(n6340), .Y(n1649) );
  OAI22XL U5899 ( .A0(n4445), .A1(n4712), .B0(n6397), .B1(n6340), .Y(n1648) );
  OAI22XL U5900 ( .A0(n4445), .A1(n4711), .B0(n6399), .B1(n6340), .Y(n1647) );
  OAI22XL U5901 ( .A0(n4445), .A1(n4710), .B0(n6401), .B1(n6340), .Y(n1646) );
  OAI22XL U5902 ( .A0(n4445), .A1(n4709), .B0(n6403), .B1(n6340), .Y(n1645) );
  OAI22XL U5903 ( .A0(n4445), .A1(n4708), .B0(n6405), .B1(n6340), .Y(n1644) );
  OAI22XL U5904 ( .A0(n4442), .A1(n4707), .B0(n6392), .B1(n6337), .Y(n1627) );
  OAI22XL U5905 ( .A0(n4442), .A1(n4706), .B0(n6394), .B1(n6337), .Y(n1626) );
  OAI22XL U5906 ( .A0(n4442), .A1(n4705), .B0(n6396), .B1(n6337), .Y(n1625) );
  OAI22XL U5907 ( .A0(n4442), .A1(n4704), .B0(n6398), .B1(n6337), .Y(n1624) );
  OAI22XL U5908 ( .A0(n4442), .A1(n4703), .B0(n6400), .B1(n6337), .Y(n1623) );
  OAI22XL U5909 ( .A0(n4442), .A1(n4702), .B0(n6402), .B1(n6337), .Y(n1622) );
  OAI22XL U5910 ( .A0(n4442), .A1(n4701), .B0(n6404), .B1(n6337), .Y(n1621) );
  OAI22XL U5911 ( .A0(n4442), .A1(n4700), .B0(n6406), .B1(n6337), .Y(n1620) );
  OAI22XL U5912 ( .A0(n4441), .A1(n4699), .B0(n6392), .B1(n6336), .Y(n1619) );
  OAI22XL U5913 ( .A0(n4441), .A1(n4698), .B0(n6394), .B1(n6336), .Y(n1618) );
  OAI22XL U5914 ( .A0(n4441), .A1(n4697), .B0(n6396), .B1(n6336), .Y(n1617) );
  OAI22XL U5915 ( .A0(n4441), .A1(n4696), .B0(n6398), .B1(n6336), .Y(n1616) );
  OAI22XL U5916 ( .A0(n4441), .A1(n4695), .B0(n6400), .B1(n6336), .Y(n1615) );
  OAI22XL U5917 ( .A0(n4441), .A1(n4694), .B0(n6402), .B1(n6336), .Y(n1614) );
  OAI22XL U5918 ( .A0(n4441), .A1(n4693), .B0(n6404), .B1(n6336), .Y(n1613) );
  OAI22XL U5919 ( .A0(n4441), .A1(n4692), .B0(n6406), .B1(n6336), .Y(n1612) );
  OAI22XL U5920 ( .A0(n4447), .A1(n4683), .B0(n6391), .B1(n6342), .Y(n1667) );
  OAI22XL U5921 ( .A0(n4447), .A1(n4682), .B0(n6393), .B1(n6342), .Y(n1666) );
  OAI22XL U5922 ( .A0(n4447), .A1(n4681), .B0(n6395), .B1(n6342), .Y(n1665) );
  OAI22XL U5923 ( .A0(n4447), .A1(n4680), .B0(n6397), .B1(n6342), .Y(n1664) );
  OAI22XL U5924 ( .A0(n4447), .A1(n4679), .B0(n6399), .B1(n6342), .Y(n1663) );
  OAI22XL U5925 ( .A0(n4447), .A1(n4678), .B0(n6401), .B1(n6342), .Y(n1662) );
  OAI22XL U5926 ( .A0(n4447), .A1(n4677), .B0(n6403), .B1(n6342), .Y(n1661) );
  OAI22XL U5927 ( .A0(n4447), .A1(n4676), .B0(n6405), .B1(n6342), .Y(n1660) );
  OAI22XL U5928 ( .A0(n4444), .A1(n4675), .B0(n6392), .B1(n6339), .Y(n1643) );
  OAI22XL U5929 ( .A0(n4444), .A1(n4674), .B0(n6394), .B1(n6339), .Y(n1642) );
  OAI22XL U5930 ( .A0(n4444), .A1(n4673), .B0(n6396), .B1(n6339), .Y(n1641) );
  OAI22XL U5931 ( .A0(n4444), .A1(n4672), .B0(n6398), .B1(n6339), .Y(n1640) );
  OAI22XL U5932 ( .A0(n4444), .A1(n4671), .B0(n6400), .B1(n6339), .Y(n1639) );
  OAI22XL U5933 ( .A0(n4444), .A1(n4670), .B0(n6402), .B1(n6339), .Y(n1638) );
  OAI22XL U5934 ( .A0(n4444), .A1(n4669), .B0(n6404), .B1(n6339), .Y(n1637) );
  OAI22XL U5935 ( .A0(n4444), .A1(n4668), .B0(n6406), .B1(n6339), .Y(n1636) );
  OAI22XL U5936 ( .A0(n4443), .A1(n4667), .B0(n6392), .B1(n6338), .Y(n1635) );
  OAI22XL U5937 ( .A0(n4443), .A1(n4666), .B0(n6394), .B1(n6338), .Y(n1634) );
  OAI22XL U5938 ( .A0(n4443), .A1(n4665), .B0(n6396), .B1(n6338), .Y(n1633) );
  OAI22XL U5939 ( .A0(n4443), .A1(n4664), .B0(n6398), .B1(n6338), .Y(n1632) );
  OAI22XL U5940 ( .A0(n4443), .A1(n4663), .B0(n6400), .B1(n6338), .Y(n1631) );
  OAI22XL U5941 ( .A0(n4443), .A1(n4662), .B0(n6402), .B1(n6338), .Y(n1630) );
  OAI22XL U5942 ( .A0(n4443), .A1(n4661), .B0(n6404), .B1(n6338), .Y(n1629) );
  OAI22XL U5943 ( .A0(n4443), .A1(n4660), .B0(n6406), .B1(n6338), .Y(n1628) );
  OAI22XL U5944 ( .A0(n4440), .A1(n4659), .B0(n6392), .B1(n6334), .Y(n1603) );
  OAI22XL U5945 ( .A0(n4440), .A1(n6046), .B0(n6394), .B1(n6334), .Y(n1602) );
  OAI22XL U5946 ( .A0(n4440), .A1(n4657), .B0(n6396), .B1(n6334), .Y(n1601) );
  OAI22XL U5947 ( .A0(n4440), .A1(n4656), .B0(n6398), .B1(n6334), .Y(n1600) );
  OAI22XL U5948 ( .A0(n4440), .A1(n4655), .B0(n6400), .B1(n6334), .Y(n1599) );
  OAI22XL U5949 ( .A0(n4440), .A1(n4654), .B0(n6402), .B1(n6334), .Y(n1598) );
  OAI22XL U5950 ( .A0(n4440), .A1(n4653), .B0(n6404), .B1(n6334), .Y(n1597) );
  OAI22XL U5951 ( .A0(n4440), .A1(n4652), .B0(n6406), .B1(n6334), .Y(n1596) );
  OAI22XL U5952 ( .A0(n4463), .A1(n4979), .B0(n6011), .B1(n6315), .Y(n1436) );
  OAI22XL U5953 ( .A0(n4463), .A1(n4984), .B0(n5980), .B1(n6315), .Y(n1432) );
  OAI22XL U5954 ( .A0(n4463), .A1(n4982), .B0(n5984), .B1(n6315), .Y(n1434) );
  OAI22XL U5955 ( .A0(n4463), .A1(n4981), .B0(n5978), .B1(n6315), .Y(n1435) );
  OAI22XL U5956 ( .A0(n4467), .A1(n4978), .B0(n6314), .B1(n4555), .Y(n1429) );
  OAI22XL U5957 ( .A0(n4451), .A1(n5033), .B0(n6003), .B1(n6310), .Y(n1319) );
  OAI22XL U5958 ( .A0(n4453), .A1(n5033), .B0(n6040), .B1(n6312), .Y(n1321) );
  OAI22XL U5959 ( .A0(n4452), .A1(n5033), .B0(n6000), .B1(n6311), .Y(n1320) );
  OAI22XL U5960 ( .A0(n4448), .A1(n4690), .B0(n6347), .B1(n4844), .Y(n1707) );
  OAI22XL U5961 ( .A0(n4448), .A1(n4689), .B0(n6394), .B1(n6347), .Y(n1706) );
  OAI22XL U5962 ( .A0(n4448), .A1(n4688), .B0(n6347), .B1(n4842), .Y(n1705) );
  OAI22XL U5963 ( .A0(n4448), .A1(n4687), .B0(n6398), .B1(n6347), .Y(n1704) );
  OAI22XL U5964 ( .A0(n4448), .A1(n4686), .B0(n6347), .B1(n4840), .Y(n1703) );
  OAI22XL U5965 ( .A0(n4448), .A1(n4685), .B0(n6347), .B1(n4838), .Y(n1701) );
  OAI22XL U5966 ( .A0(n4448), .A1(n4684), .B0(n6347), .B1(n4837), .Y(n1700) );
  OA21XL U5967 ( .A0(\add_653_S2/carry[3] ), .A1(n6313), .B0(n5006), .Y(n4920)
         );
  CLKBUFX3 U5968 ( .A(n4936), .Y(n6341) );
  NAND2X1 U5969 ( .A(n4934), .B(n4929), .Y(n4936) );
  CLKBUFX3 U5970 ( .A(n4935), .Y(n6342) );
  NAND2X1 U5971 ( .A(n4934), .B(n4927), .Y(n4935) );
  CLKBUFX3 U5972 ( .A(n4965), .Y(n6319) );
  NAND2X1 U5973 ( .A(n4966), .B(n4924), .Y(n4965) );
  CLKBUFX3 U5974 ( .A(n4967), .Y(n6318) );
  NAND2X1 U5975 ( .A(n4966), .B(n4927), .Y(n4967) );
  CLKBUFX3 U5976 ( .A(n4952), .Y(n6329) );
  NAND2X1 U5977 ( .A(n4950), .B(n4929), .Y(n4952) );
  CLKBUFX3 U5978 ( .A(n4953), .Y(n6328) );
  NAND2X1 U5979 ( .A(n4950), .B(n4931), .Y(n4953) );
  CLKBUFX3 U5980 ( .A(n4958), .Y(n6325) );
  NAND2X1 U5981 ( .A(n4956), .B(n4929), .Y(n4958) );
  CLKBUFX3 U5982 ( .A(n4959), .Y(n6324) );
  NAND2X1 U5983 ( .A(n4956), .B(n4931), .Y(n4959) );
  CLKBUFX3 U5984 ( .A(n4963), .Y(n6321) );
  NAND2X1 U5985 ( .A(n4961), .B(n4929), .Y(n4963) );
  CLKBUFX3 U5986 ( .A(n4964), .Y(n6320) );
  NAND2X1 U5987 ( .A(n4961), .B(n4931), .Y(n4964) );
  CLKBUFX3 U5988 ( .A(n4949), .Y(n6331) );
  NAND2X1 U5989 ( .A(n4950), .B(n4924), .Y(n4949) );
  CLKBUFX3 U5990 ( .A(n4955), .Y(n6327) );
  NAND2X1 U5991 ( .A(n4956), .B(n4924), .Y(n4955) );
  CLKBUFX3 U5992 ( .A(n4957), .Y(n6326) );
  NAND2X1 U5993 ( .A(n4956), .B(n4927), .Y(n4957) );
  CLKBUFX3 U5994 ( .A(n4960), .Y(n6323) );
  NAND2X1 U5995 ( .A(n4961), .B(n4924), .Y(n4960) );
  CLKBUFX3 U5996 ( .A(n4962), .Y(n6322) );
  NAND2X1 U5997 ( .A(n4961), .B(n4927), .Y(n4962) );
  CLKBUFX3 U5998 ( .A(n4941), .Y(n6337) );
  NAND2X1 U5999 ( .A(n4939), .B(n4929), .Y(n4941) );
  CLKBUFX3 U6000 ( .A(n4942), .Y(n6336) );
  NAND2X1 U6001 ( .A(n4939), .B(n4931), .Y(n4942) );
  CLKBUFX3 U6002 ( .A(n4938), .Y(n6339) );
  NAND2X1 U6003 ( .A(n4939), .B(n4924), .Y(n4938) );
  CLKBUFX3 U6004 ( .A(n4940), .Y(n6338) );
  NAND2X1 U6005 ( .A(n4939), .B(n4927), .Y(n4940) );
  CLKBUFX3 U6006 ( .A(n4945), .Y(n6334) );
  NAND2X1 U6007 ( .A(n4944), .B(n4927), .Y(n4945) );
  CLKBUFX3 U6008 ( .A(n4937), .Y(n6340) );
  NAND2X1 U6009 ( .A(n4934), .B(n4931), .Y(n4937) );
  CLKBUFX3 U6010 ( .A(n4923), .Y(n6347) );
  NAND2X1 U6011 ( .A(n4924), .B(n4925), .Y(n4923) );
  OAI222XL U6012 ( .A0(n6361), .A1(n4669), .B0(n6368), .B1(n4733), .C0(n6352), 
        .C1(n4757), .Y(n5707) );
  OAI222XL U6013 ( .A0(n6360), .A1(n4674), .B0(n6368), .B1(n4738), .C0(n6352), 
        .C1(n6012), .Y(n5711) );
  OAI222XL U6014 ( .A0(n6357), .A1(n4672), .B0(n6368), .B1(n4736), .C0(n6352), 
        .C1(n4760), .Y(n5715) );
  OAI222X1 U6015 ( .A0(n4617), .A1(n5403), .B0(n5374), .B1(n5404), .C0(n5405), 
        .C1(n5984), .Y(n5359) );
  OAI222X1 U6016 ( .A0(n4619), .A1(n5403), .B0(n5369), .B1(n5404), .C0(n5405), 
        .C1(n6011), .Y(n5363) );
  OAI31X1 U6017 ( .A0(n5071), .A1(n4858), .A2(n5072), .B0(n5073), .Y(n5045) );
  OAI221XL U6018 ( .A0(n5074), .A1(n5075), .B0(n4507), .B1(n5076), .C0(n4858), 
        .Y(n5073) );
  AO22X1 U6019 ( .A0(n5077), .A1(n4542), .B0(n5078), .B1(n4548), .Y(n5072) );
  OAI222XL U6020 ( .A0(n4510), .A1(n5080), .B0(n5081), .B1(n5075), .C0(n4508), 
        .C1(n5070), .Y(n5071) );
  NAND4BX1 U6021 ( .AN(n5141), .B(n4830), .C(n5142), .D(n5143), .Y(n5140) );
  OAI21X2 U6022 ( .A0(n4911), .A1(n4458), .B0(n4845), .Y(n4922) );
  OAI222XL U6023 ( .A0(n6357), .A1(n4668), .B0(n6368), .B1(n4732), .C0(n6352), 
        .C1(n4756), .Y(n5719) );
  OAI222XL U6024 ( .A0(n6357), .A1(n4675), .B0(n6368), .B1(n4739), .C0(n6352), 
        .C1(n4763), .Y(n5722) );
  NAND4X1 U6025 ( .A(n5277), .B(n5278), .C(n5279), .D(n5280), .Y(n5084) );
  XNOR2X1 U6026 ( .A(n5255), .B(n5201), .Y(n5278) );
  XOR2X1 U6027 ( .A(n5257), .B(n5205), .Y(n5277) );
  NOR4X1 U6028 ( .A(n5281), .B(n5282), .C(n5283), .D(n5284), .Y(n5280) );
  NAND4X1 U6029 ( .A(n5301), .B(n5302), .C(n5303), .D(n5304), .Y(n5085) );
  XOR2X1 U6030 ( .A(n5248), .B(n5243), .Y(n5301) );
  XOR2X1 U6031 ( .A(n5246), .B(n5241), .Y(n5302) );
  NOR4X1 U6032 ( .A(n5305), .B(n5306), .C(n5307), .D(n5308), .Y(n5304) );
  XOR2X1 U6033 ( .A(n5355), .B(n5416), .Y(n5415) );
  AOI32X1 U6034 ( .A0(n6348), .A1(n6021), .A2(n4609), .B0(n5103), .B1(n5104), 
        .Y(n5099) );
  NOR4X1 U6035 ( .A(n5112), .B(n5113), .C(n5114), .D(n5115), .Y(n5103) );
  XOR2X1 U6036 ( .A(n5117), .B(n4591), .Y(n5114) );
  NAND4X1 U6037 ( .A(n5264), .B(n5265), .C(n5266), .D(n5267), .Y(n5102) );
  XOR2X1 U6038 ( .A(n5342), .B(n5185), .Y(n5265) );
  XNOR2X1 U6039 ( .A(n5173), .B(n5254), .Y(n5264) );
  NOR4X1 U6040 ( .A(n5268), .B(n5269), .C(n5270), .D(n5271), .Y(n5267) );
  OAI22XL U6041 ( .A0(n5079), .A1(n5084), .B0(n5085), .B1(n5070), .Y(n5083) );
  OAI22XL U6042 ( .A0(n4834), .A1(n4912), .B0(n4859), .B1(n4913), .Y(n1450) );
  OAI22XL U6043 ( .A0(n4860), .A1(n4912), .B0(n4858), .B1(n4913), .Y(n1722) );
  OAI22XL U6044 ( .A0(n4834), .A1(n4972), .B0(n4973), .B1(n4846), .Y(n1448) );
  XOR2X1 U6045 ( .A(n5191), .B(n4586), .Y(n5275) );
  XOR2X1 U6046 ( .A(n5256), .B(n5165), .Y(n5276) );
  XOR2X1 U6047 ( .A(n5203), .B(n4583), .Y(n5287) );
  XOR2X1 U6048 ( .A(n5200), .B(n4590), .Y(n5288) );
  XOR2X1 U6049 ( .A(n5249), .B(n4563), .Y(n5299) );
  XOR2X1 U6050 ( .A(n5219), .B(n4569), .Y(n5300) );
  XNOR2X1 U6051 ( .A(n5375), .B(n5358), .Y(n5406) );
  OAI21XL U6052 ( .A0(n4457), .A1(n4857), .B0(n4912), .Y(n1449) );
  CLKBUFX3 U6053 ( .A(n4843), .Y(n6393) );
  CLKBUFX3 U6054 ( .A(n4930), .Y(n6344) );
  NAND2X1 U6055 ( .A(n4931), .B(n4925), .Y(n4930) );
  CLKBUFX3 U6056 ( .A(n4928), .Y(n6345) );
  NAND2X1 U6057 ( .A(n4929), .B(n4925), .Y(n4928) );
  CLKBUFX3 U6058 ( .A(n4926), .Y(n6346) );
  NAND2X1 U6059 ( .A(n4927), .B(n4925), .Y(n4926) );
  CLKBUFX3 U6060 ( .A(n4968), .Y(n6317) );
  NAND2X1 U6061 ( .A(n4966), .B(n4929), .Y(n4968) );
  CLKBUFX3 U6062 ( .A(n4951), .Y(n6330) );
  NAND2X1 U6063 ( .A(n4950), .B(n4927), .Y(n4951) );
  CLKBUFX3 U6064 ( .A(n4946), .Y(n6333) );
  NAND2X1 U6065 ( .A(n4944), .B(n4929), .Y(n4946) );
  CLKBUFX3 U6066 ( .A(n4943), .Y(n6335) );
  NAND2X1 U6067 ( .A(n4944), .B(n4924), .Y(n4943) );
  CLKBUFX3 U6068 ( .A(n4933), .Y(n6343) );
  NAND2X1 U6069 ( .A(n4934), .B(n4924), .Y(n4933) );
  AO21X1 U6070 ( .A0(n5011), .A1(n5067), .B0(n4849), .Y(n5066) );
  OAI222X1 U6071 ( .A0(n6353), .A1(n4735), .B0(n6361), .B1(n4759), .C0(n6371), 
        .C1(n4671), .Y(n5581) );
  OAI222X1 U6072 ( .A0(n6353), .A1(n4739), .B0(n6361), .B1(n4763), .C0(n6371), 
        .C1(n4675), .Y(n5585) );
  OAI222X1 U6073 ( .A0(n6353), .A1(n4732), .B0(n6362), .B1(n4756), .C0(n6371), 
        .C1(n4668), .Y(n5648) );
  OAI222X1 U6074 ( .A0(n6353), .A1(n4736), .B0(n6361), .B1(n4760), .C0(n6371), 
        .C1(n4672), .Y(n5814) );
  OAI222X1 U6075 ( .A0(n6353), .A1(n4738), .B0(n6361), .B1(n6012), .C0(n6371), 
        .C1(n4674), .Y(n5775) );
  OAI222X1 U6076 ( .A0(n6353), .A1(n4733), .B0(n6361), .B1(n4757), .C0(n6371), 
        .C1(n4669), .Y(n5651) );
  OAI222X1 U6077 ( .A0(n6353), .A1(n4737), .B0(n6361), .B1(n4761), .C0(n6371), 
        .C1(n4673), .Y(n5828) );
  OAI222X1 U6078 ( .A0(n6353), .A1(n4734), .B0(n6361), .B1(n4758), .C0(n6371), 
        .C1(n4670), .Y(n5820) );
  OAI222X1 U6079 ( .A0(n5561), .A1(n6387), .B0(n5623), .B1(n6385), .C0(
        match_index[1]), .C1(n4636), .Y(n5653) );
  OAI222X1 U6080 ( .A0(n5850), .A1(n6387), .B0(n5779), .B1(n6386), .C0(
        match_index[1]), .C1(n4618), .Y(n5813) );
  OAI222X1 U6081 ( .A0(n6387), .A1(n5651), .B0(n4630), .B1(n6386), .C0(
        match_index[1]), .C1(n4631), .Y(n5673) );
  OAI222X1 U6082 ( .A0(n5357), .A1(n5403), .B0(n5381), .B1(n5404), .C0(n5405), 
        .C1(n5980), .Y(n5356) );
  OAI222X1 U6083 ( .A0(n4612), .A1(n5403), .B0(n5375), .B1(n5404), .C0(n5405), 
        .C1(n5978), .Y(n5358) );
  AOI222XL U6084 ( .A0(n4474), .A1(n4475), .B0(n5464), .B1(n4478), .C0(n5436), 
        .C1(n5465), .Y(n5463) );
  CLKINVX1 U6085 ( .A(n5469), .Y(n4474) );
  CLKINVX1 U6086 ( .A(n5468), .Y(n4478) );
  NAND2X2 U6087 ( .A(n5405), .B(n5403), .Y(n5404) );
  AOI221XL U6088 ( .A0(n4828), .A1(n5078), .B0(n4829), .B1(n5082), .C0(n5128), 
        .Y(n5096) );
  CLKINVX1 U6089 ( .A(n4974), .Y(n4828) );
  OAI32X1 U6090 ( .A0(n4509), .A1(n6348), .A2(n4834), .B0(n4510), .B1(n4973), 
        .Y(n5128) );
  CLKINVX1 U6091 ( .A(n5077), .Y(n4509) );
  OAI22XL U6092 ( .A0(n6013), .A1(n5694), .B0(n4640), .B1(n5695), .Y(n5693) );
  OA22X1 U6093 ( .A0(n6457), .A1(n5682), .B0(n6296), .B1(n5709), .Y(n5369) );
  OA22X1 U6094 ( .A0(n6457), .A1(n5778), .B0(n6296), .B1(n5713), .Y(n5374) );
  OA22X1 U6095 ( .A0(n6457), .A1(n5782), .B0(n6297), .B1(n5725), .Y(n5381) );
  OAI22XL U6096 ( .A0(n5985), .A1(n5694), .B0(n4610), .B1(n5695), .Y(n5704) );
  OAI22XL U6097 ( .A0(n6033), .A1(n5694), .B0(n4619), .B1(n5695), .Y(n5708) );
  OAI22XL U6098 ( .A0(n6034), .A1(n5694), .B0(n4617), .B1(n5695), .Y(n5712) );
  AOI222XL U6099 ( .A0(n5698), .A1(n5735), .B0(n4628), .B1(n5700), .C0(n4623), 
        .C1(n5701), .Y(n5734) );
  OAI222XL U6100 ( .A0(n6361), .A1(n4673), .B0(n6368), .B1(n4737), .C0(n6352), 
        .C1(n4761), .Y(n5735) );
  NAND2X2 U6101 ( .A(n5405), .B(n5149), .Y(n5403) );
  NAND4X1 U6102 ( .A(n5224), .B(n5225), .C(n5226), .D(n5227), .Y(n5136) );
  NOR4X1 U6103 ( .A(n5228), .B(n5229), .C(n5230), .D(n5231), .Y(n5227) );
  NAND4X1 U6104 ( .A(n5175), .B(n5176), .C(n5177), .D(n5178), .Y(n5138) );
  XOR2X1 U6105 ( .A(n5257), .B(n5258), .Y(n5175) );
  XNOR2X1 U6106 ( .A(n5255), .B(n5256), .Y(n5176) );
  NOR4X1 U6107 ( .A(n5179), .B(n5180), .C(n5181), .D(n5182), .Y(n5178) );
  NAND4X1 U6108 ( .A(n5209), .B(n5210), .C(n5211), .D(n5212), .Y(n5132) );
  XOR2X1 U6109 ( .A(n5248), .B(n5249), .Y(n5209) );
  XOR2X1 U6110 ( .A(n5246), .B(n5247), .Y(n5210) );
  NOR4X1 U6111 ( .A(n5213), .B(n5214), .C(n5215), .D(n5216), .Y(n5212) );
  NOR3X1 U6112 ( .A(n5676), .B(n5442), .C(n5677), .Y(n5665) );
  OAI22XL U6113 ( .A0(n4585), .A1(n5679), .B0(n6035), .B1(n5680), .Y(n5812) );
  OAI21XL U6114 ( .A0(n5441), .A1(n5442), .B0(n5443), .Y(n5439) );
  NAND4X1 U6115 ( .A(n5436), .B(n4595), .C(n4591), .D(n5923), .Y(n5430) );
  NAND4BX1 U6116 ( .AN(n5435), .B(n5450), .C(n5451), .D(n5386), .Y(n5433) );
  NOR3X1 U6117 ( .A(n5594), .B(n5449), .C(n5595), .Y(n5565) );
  XOR2X1 U6118 ( .A(n5884), .B(n5885), .Y(n5594) );
  XNOR2X1 U6119 ( .A(n5255), .B(n5596), .Y(n5595) );
  OAI22XL U6120 ( .A0(n4583), .A1(n5597), .B0(n6053), .B1(n5598), .Y(n5885) );
  NOR3X1 U6121 ( .A(n5630), .B(n5448), .C(n5631), .Y(n5605) );
  XNOR2X1 U6122 ( .A(n5251), .B(n5862), .Y(n5630) );
  XOR2X1 U6123 ( .A(n5632), .B(n5633), .Y(n5631) );
  OAI22XL U6124 ( .A0(n5251), .A1(n5634), .B0(n6058), .B1(n5863), .Y(n5862) );
  NOR3X1 U6125 ( .A(n5661), .B(n5662), .C(n5445), .Y(n5639) );
  XOR2X1 U6126 ( .A(n5832), .B(n4575), .Y(n5662) );
  XOR2X1 U6127 ( .A(n5840), .B(n5841), .Y(n5661) );
  OAI22XL U6128 ( .A0(n4492), .A1(n6049), .B0(n5337), .B1(n5833), .Y(n5832) );
  NOR3X1 U6129 ( .A(n5235), .B(n5236), .C(n5237), .Y(n5226) );
  NOR3X1 U6130 ( .A(n5189), .B(n5134), .C(n5190), .Y(n5177) );
  XOR2X1 U6131 ( .A(n5254), .B(n4583), .Y(n5189) );
  XOR2X1 U6132 ( .A(n5191), .B(n4590), .Y(n5190) );
  NOR3X1 U6133 ( .A(n5206), .B(n5132), .C(n5207), .Y(n5194) );
  XOR2X1 U6134 ( .A(n5250), .B(n4563), .Y(n5206) );
  XOR2X1 U6135 ( .A(n5208), .B(n4569), .Y(n5207) );
  NAND2X1 U6136 ( .A(n5048), .B(n4471), .Y(n5043) );
  NAND4X1 U6137 ( .A(n5049), .B(n5050), .C(n5051), .D(n5052), .Y(n5048) );
  XOR2X1 U6138 ( .A(n6476), .B(N247), .Y(n5050) );
  AOI2BB2X1 U6139 ( .B0(n5436), .B1(n5437), .A0N(n5438), .A1N(n5436), .Y(n5434) );
  OAI22XL U6140 ( .A0(n5446), .A1(n4551), .B0(n5447), .B1(n5444), .Y(n5437) );
  AOI221XL U6141 ( .A0(n4537), .A1(n4546), .B0(n4545), .B1(n5439), .C0(n5440), 
        .Y(n5438) );
  OA21XL U6142 ( .A0(n5056), .A1(n5448), .B0(n5449), .Y(n5446) );
  NAND4BX1 U6143 ( .AN(n5457), .B(n5458), .C(n5459), .D(n5460), .Y(n5432) );
  OAI21XL U6144 ( .A0(n4506), .A1(n5454), .B0(n5461), .Y(n5460) );
  NAND3X1 U6145 ( .A(n5470), .B(n6349), .C(n4514), .Y(n5458) );
  OAI2BB1X1 U6146 ( .A0N(n5480), .A1N(match_index[4]), .B0(n5387), .Y(n5457)
         );
  NOR3X1 U6147 ( .A(n5260), .B(n5169), .C(n5168), .Y(n5496) );
  NOR2X1 U6148 ( .A(n5449), .B(n5056), .Y(n5464) );
  NAND3X1 U6149 ( .A(n4475), .B(n5550), .C(n5551), .Y(n5533) );
  OAI21XL U6150 ( .A0(n4565), .A1(n6052), .B0(n5556), .Y(n5550) );
  XOR2X1 U6151 ( .A(n5552), .B(n5165), .Y(n5551) );
  OAI21XL U6152 ( .A0(n4565), .A1(n4473), .B0(n6052), .Y(n5556) );
  CLKBUFX3 U6153 ( .A(n451), .Y(n6477) );
  CLKBUFX3 U6154 ( .A(n6461), .Y(n6464) );
  CLKBUFX3 U6155 ( .A(n6461), .Y(n6463) );
  CLKBUFX3 U6156 ( .A(n6460), .Y(n6454) );
  CLKINVX1 U6157 ( .A(n6451), .Y(n6460) );
  CLKBUFX3 U6158 ( .A(n6469), .Y(n6467) );
  CLKBUFX3 U6159 ( .A(n6469), .Y(n6468) );
  CLKBUFX3 U6160 ( .A(n6469), .Y(n6466) );
  OAI222X1 U6161 ( .A0(n6384), .A1(n5822), .B0(n4603), .B1(n6381), .C0(n453), 
        .C1(n5512), .Y(n5542) );
  CLKINVX1 U6162 ( .A(n5513), .Y(n4603) );
  OAI221XL U6163 ( .A0(n5600), .A1(n6385), .B0(n6382), .B1(n5775), .C0(n5878), 
        .Y(n5857) );
  OAI221XL U6164 ( .A0(n5357), .A1(n5695), .B0(n6014), .B1(n5694), .C0(n5724), 
        .Y(n5723) );
  XOR2X1 U6165 ( .A(n5239), .B(n4598), .Y(n5308) );
  XOR2X1 U6166 ( .A(n5218), .B(n4589), .Y(n5296) );
  XOR2X1 U6167 ( .A(n5233), .B(n4588), .Y(n5307) );
  XOR2X1 U6168 ( .A(n5217), .B(n4599), .Y(n5293) );
  XOR2X1 U6169 ( .A(n5238), .B(n4568), .Y(n5306) );
  OAI22XL U6170 ( .A0(n4612), .A1(n5695), .B0(n6032), .B1(n5694), .Y(n5729) );
  OAI22XL U6171 ( .A0(n4581), .A1(n5679), .B0(n5992), .B1(n5680), .Y(n5678) );
  OA22X1 U6172 ( .A0(n4868), .A1(n5310), .B0(n4584), .B1(n5309), .Y(n5241) );
  CLKINVX1 U6173 ( .A(n5338), .Y(n4576) );
  OAI221XL U6174 ( .A0(n4867), .A1(n5310), .B0(n5309), .B1(n5337), .C0(n5135), 
        .Y(n5338) );
  CLKINVX1 U6175 ( .A(n5376), .Y(n4554) );
  OA22X1 U6176 ( .A0(n5986), .A1(n5298), .B0(n5204), .B1(n5297), .Y(n5247) );
  OA22X1 U6177 ( .A0(n6051), .A1(n5298), .B0(n5251), .B1(n5297), .Y(n5245) );
  OA22X1 U6178 ( .A0(n4869), .A1(n5310), .B0(n4593), .B1(n5309), .Y(n5232) );
  OA22X1 U6179 ( .A0(n4870), .A1(n5310), .B0(n5221), .B1(n5309), .Y(n5234) );
  OA22X1 U6180 ( .A0(n6023), .A1(n5298), .B0(n5202), .B1(n5297), .Y(n5220) );
  CLKBUFX3 U6181 ( .A(n4844), .Y(n6391) );
  CLKBUFX3 U6182 ( .A(n4842), .Y(n6395) );
  CLKBUFX3 U6183 ( .A(n4841), .Y(n6397) );
  CLKBUFX3 U6184 ( .A(n4840), .Y(n6399) );
  CLKBUFX3 U6185 ( .A(n4839), .Y(n6401) );
  CLKBUFX3 U6186 ( .A(n4838), .Y(n6403) );
  CLKBUFX3 U6187 ( .A(n4837), .Y(n6405) );
  CLKBUFX3 U6188 ( .A(n6461), .Y(n6465) );
  CLKBUFX3 U6189 ( .A(n451), .Y(n6476) );
  CLKINVX1 U6190 ( .A(n6453), .Y(n6459) );
  CLKINVX1 U6191 ( .A(n5508), .Y(n4602) );
  CLKINVX1 U6192 ( .A(n5593), .Y(n4607) );
  CLKINVX1 U6193 ( .A(n5503), .Y(n4601) );
  CLKINVX1 U6194 ( .A(n5872), .Y(n4605) );
  CLKINVX1 U6195 ( .A(n5866), .Y(n4606) );
  CLKINVX1 U6196 ( .A(n5602), .Y(n4604) );
  OAI211X1 U6197 ( .A0(n5931), .A1(n6388), .B0(n5526), .C0(n5932), .Y(n5521)
         );
  AOI222XL U6198 ( .A0(match_index[3]), .A1(n4740), .B0(n6376), .B1(n4652), 
        .C0(match_index[4]), .C1(n4812), .Y(n5931) );
  OA22X1 U6199 ( .A0(n6385), .A1(n5620), .B0(match_index[1]), .B1(n5621), .Y(
        n5932) );
  OAI211X1 U6200 ( .A0(n5543), .A1(n6388), .B0(n5526), .C0(n5544), .Y(n5510)
         );
  AOI222XL U6201 ( .A0(match_index[3]), .A1(n4742), .B0(n6376), .B1(n4654), 
        .C0(match_index[4]), .C1(n4814), .Y(n5543) );
  OA22X1 U6202 ( .A0(n6385), .A1(n5545), .B0(match_index[1]), .B1(n5546), .Y(
        n5544) );
  OAI211X1 U6203 ( .A0(n5559), .A1(n6388), .B0(n5526), .C0(n5560), .Y(n5499)
         );
  AOI222XL U6204 ( .A0(match_index[3]), .A1(n4747), .B0(n6378), .B1(n4659), 
        .C0(match_index[4]), .C1(n4819), .Y(n5559) );
  OA22X1 U6205 ( .A0(n6386), .A1(n5561), .B0(match_index[1]), .B1(n5562), .Y(
        n5560) );
  OAI211X1 U6206 ( .A0(n5524), .A1(n6388), .B0(n5526), .C0(n5527), .Y(n5505)
         );
  AOI222XL U6207 ( .A0(match_index[3]), .A1(n4743), .B0(n6376), .B1(n4655), 
        .C0(match_index[4]), .C1(n4815), .Y(n5524) );
  OA22X1 U6208 ( .A0(n6386), .A1(n5529), .B0(match_index[1]), .B1(n5530), .Y(
        n5527) );
  OAI211X1 U6209 ( .A0(n5953), .A1(n6388), .B0(n5526), .C0(n5954), .Y(n5532)
         );
  AOI222XL U6210 ( .A0(match_index[3]), .A1(n4741), .B0(n6375), .B1(n4653), 
        .C0(match_index[4]), .C1(n4813), .Y(n5953) );
  OA22X1 U6211 ( .A0(n6385), .A1(n5616), .B0(match_index[1]), .B1(n5617), .Y(
        n5954) );
  OAI211X1 U6212 ( .A0(n5943), .A1(n6388), .B0(n5526), .C0(n5944), .Y(n5549)
         );
  AOI222XL U6213 ( .A0(match_index[3]), .A1(n4745), .B0(n6376), .B1(n4657), 
        .C0(match_index[4]), .C1(n4817), .Y(n5943) );
  OA22X1 U6214 ( .A0(n6385), .A1(n5844), .B0(match_index[1]), .B1(n5892), .Y(
        n5944) );
  NAND4BX1 U6215 ( .AN(n5386), .B(n5387), .C(n4514), .D(n5388), .Y(n5067) );
  NOR3X1 U6216 ( .A(n5389), .B(n5390), .C(n5391), .Y(n5388) );
  XOR2X1 U6217 ( .A(match_index[4]), .B(n5394), .Y(n5389) );
  XOR2X1 U6218 ( .A(n5217), .B(n4598), .Y(n5216) );
  XOR2X1 U6219 ( .A(n5200), .B(n4589), .Y(n5199) );
  XOR2X1 U6220 ( .A(n5118), .B(n4565), .Y(n5163) );
  XOR2X1 U6221 ( .A(n5116), .B(n4572), .Y(n5115) );
  XOR2X1 U6222 ( .A(n5218), .B(n4588), .Y(n5215) );
  XOR2X1 U6223 ( .A(n5108), .B(n4595), .Y(n5107) );
  XOR2X1 U6224 ( .A(n5250), .B(n4564), .Y(n5283) );
  XOR2X1 U6225 ( .A(n5185), .B(n4564), .Y(n5181) );
  XOR2X1 U6226 ( .A(n5208), .B(n4570), .Y(n5281) );
  XOR2X1 U6227 ( .A(n5188), .B(n4570), .Y(n5179) );
  XOR2X1 U6228 ( .A(n5205), .B(n4599), .Y(n5196) );
  XOR2X1 U6229 ( .A(n5118), .B(n4566), .Y(n5113) );
  XOR2X1 U6230 ( .A(n5258), .B(n4596), .Y(n5270) );
  XOR2X1 U6231 ( .A(n5219), .B(n4568), .Y(n5214) );
  XOR2X1 U6232 ( .A(n5188), .B(n4571), .Y(n5269) );
  OAI22XL U6233 ( .A0(n4490), .A1(n6057), .B0(n4574), .B1(n5634), .Y(n5633) );
  NOR4X1 U6234 ( .A(n5161), .B(n5162), .C(n5163), .D(n5164), .Y(n5160) );
  XOR2X1 U6235 ( .A(n5122), .B(n5165), .Y(n5164) );
  XOR2X1 U6236 ( .A(n5116), .B(n4571), .Y(n5162) );
  NAND2X1 U6237 ( .A(n5170), .B(n5171), .Y(n5161) );
  OAI22XL U6238 ( .A0(n4538), .A1(n6041), .B0(n4577), .B1(n5679), .Y(n5818) );
  OAI22XL U6239 ( .A0(n4593), .A1(n5833), .B0(n6050), .B1(n5842), .Y(n5841) );
  OAI22XL U6240 ( .A0(n4594), .A1(n5679), .B0(n6042), .B1(n5680), .Y(n5824) );
  OAI22XL U6241 ( .A0(n5204), .A1(n5634), .B0(n6043), .B1(n5863), .Y(n5869) );
  OAI22XL U6242 ( .A0(n5221), .A1(n5833), .B0(n5994), .B1(n5842), .Y(n5854) );
  OAI22XL U6243 ( .A0(n4584), .A1(n5833), .B0(n6036), .B1(n5842), .Y(n5848) );
  NAND2X1 U6244 ( .A(n5135), .B(n5309), .Y(n5310) );
  NAND3X1 U6245 ( .A(n6025), .B(n5987), .C(n5343), .Y(n5137) );
  NAND3X1 U6246 ( .A(n6024), .B(n5988), .C(n5341), .Y(n5133) );
  NAND3X1 U6247 ( .A(n6026), .B(n5989), .C(n5263), .Y(n5155) );
  NAND3X1 U6248 ( .A(n6023), .B(n5986), .C(n5340), .Y(n5130) );
  NAND3X1 U6249 ( .A(n4870), .B(n4868), .C(n5339), .Y(n5135) );
  CLKINVX1 U6250 ( .A(n5168), .Y(n4566) );
  CLKINVX1 U6251 ( .A(n5169), .Y(n4572) );
  CLKINVX1 U6252 ( .A(n5260), .Y(n4579) );
  NAND2X1 U6253 ( .A(n5376), .B(n5345), .Y(n5371) );
  CLKINVX1 U6254 ( .A(n5121), .Y(n4580) );
  CLKINVX1 U6255 ( .A(n5123), .Y(n4582) );
  NAND3X1 U6256 ( .A(n4878), .B(n4876), .C(n5385), .Y(n5345) );
  NAND2X1 U6257 ( .A(n4516), .B(n4857), .Y(n5472) );
  CLKINVX1 U6258 ( .A(n5259), .Y(n4505) );
  OAI221XL U6259 ( .A0(n6063), .A1(n5166), .B0(n4579), .B1(n5167), .C0(n5155), 
        .Y(n5259) );
  OA22X1 U6260 ( .A0(n5989), .A1(n5166), .B0(n4582), .B1(n5167), .Y(n5124) );
  OA22X1 U6261 ( .A0(n6070), .A1(n5166), .B0(n4591), .B1(n5167), .Y(n5117) );
  OA22X1 U6262 ( .A0(n6026), .A1(n5166), .B0(n4580), .B1(n5167), .Y(n5122) );
  OA22X1 U6263 ( .A0(n6024), .A1(n5285), .B0(n5255), .B1(n5286), .Y(n5201) );
  OA22X1 U6264 ( .A0(n6059), .A1(n5285), .B0(n5187), .B1(n5286), .Y(n5252) );
  OA22X1 U6265 ( .A0(n5987), .A1(n5273), .B0(n5173), .B1(n5274), .Y(n5254) );
  OA22X1 U6266 ( .A0(n6025), .A1(n5273), .B0(n5165), .B1(n5274), .Y(n5256) );
  OA22X1 U6267 ( .A0(n5988), .A1(n5285), .B0(n4583), .B1(n5286), .Y(n5203) );
  OA22X1 U6268 ( .A0(n6065), .A1(n5273), .B0(n4592), .B1(n5274), .Y(n5186) );
  CLKINVX1 U6269 ( .A(n5475), .Y(n4512) );
  NAND2X1 U6270 ( .A(n5119), .B(n5120), .Y(n5112) );
  XOR2X1 U6271 ( .A(n5121), .B(n5122), .Y(n5120) );
  XOR2X1 U6272 ( .A(n5123), .B(n5124), .Y(n5119) );
  OAI211X1 U6273 ( .A0(n5918), .A1(n6388), .B0(n5526), .C0(n5919), .Y(n5539)
         );
  AOI222XL U6274 ( .A0(match_index[3]), .A1(n4744), .B0(n6376), .B1(n4656), 
        .C0(match_index[4]), .C1(n4816), .Y(n5918) );
  OA22X1 U6275 ( .A0(n6385), .A1(n5850), .B0(match_index[1]), .B1(n5886), .Y(
        n5919) );
  OAI211X1 U6276 ( .A0(n5909), .A1(n6388), .B0(n5526), .C0(n5910), .Y(n5554)
         );
  AOI222XL U6277 ( .A0(match_index[3]), .A1(n4746), .B0(n6376), .B1(n6046), 
        .C0(match_index[4]), .C1(n4818), .Y(n5909) );
  OA22X1 U6278 ( .A0(n6386), .A1(n5858), .B0(match_index[1]), .B1(n5882), .Y(
        n5910) );
  XOR2X1 U6279 ( .A(n5272), .B(n5541), .Y(n5535) );
  OAI22XL U6280 ( .A0(n4473), .A1(n6068), .B0(n4578), .B1(n5520), .Y(n5541) );
  XNOR2X1 U6281 ( .A(n5173), .B(n5537), .Y(n5536) );
  OAI22XL U6282 ( .A0(n5173), .A1(n5520), .B0(n6005), .B1(n5538), .Y(n5537) );
  XOR2X1 U6283 ( .A(n5172), .B(n5547), .Y(n5534) );
  OAI22XL U6284 ( .A0(n4592), .A1(n5520), .B0(n6069), .B1(n5538), .Y(n5547) );
  NAND2X1 U6285 ( .A(n5462), .B(n5679), .Y(n5680) );
  XOR2X1 U6286 ( .A(n5261), .B(n5110), .Y(n5158) );
  OAI22XL U6287 ( .A0(n4477), .A1(n6062), .B0(n4573), .B1(n5597), .Y(n5896) );
  OAI22XL U6288 ( .A0(n5255), .A1(n5597), .B0(n6001), .B1(n5598), .Y(n5596) );
  OAI22XL U6289 ( .A0(n5165), .A1(n5520), .B0(n6060), .B1(n5538), .Y(n5552) );
  OAI22XL U6290 ( .A0(n5187), .A1(n5597), .B0(n6064), .B1(n5598), .Y(n5890) );
  OAI22XL U6291 ( .A0(n5202), .A1(n5634), .B0(n5998), .B1(n5863), .Y(n5875) );
  NAND2X1 U6292 ( .A(n5130), .B(n5297), .Y(n5298) );
  NAND2X1 U6293 ( .A(n5133), .B(n5286), .Y(n5285) );
  CLKINVX1 U6294 ( .A(n5461), .Y(n4514) );
  OAI21XL U6295 ( .A0(n4471), .A1(n5016), .B0(n5011), .Y(N842) );
  CLKINVX1 U6296 ( .A(n5679), .Y(n4538) );
  NAND3X1 U6297 ( .A(n5992), .B(n6035), .C(n5825), .Y(n5462) );
  AND4X1 U6298 ( .A(n5111), .B(n5435), .C(n4551), .D(n4545), .Y(n5923) );
  NAND2X1 U6299 ( .A(n5468), .B(n5597), .Y(n5598) );
  NAND2X1 U6300 ( .A(n5467), .B(n5634), .Y(n5863) );
  NAND2X1 U6301 ( .A(n5466), .B(n5833), .Y(n5842) );
  NAND2X1 U6302 ( .A(n5137), .B(n5274), .Y(n5273) );
  NAND2X1 U6303 ( .A(n5155), .B(n5167), .Y(n5166) );
  CLKINVX1 U6304 ( .A(n5394), .Y(n4506) );
  CLKINVX1 U6305 ( .A(N166), .Y(n4833) );
  NAND4X1 U6306 ( .A(n5996), .B(n5979), .C(n6037), .D(n5981), .Y(n5740) );
  NAND3X1 U6307 ( .A(n5994), .B(n6036), .C(n5855), .Y(n5466) );
  CLKINVX1 U6308 ( .A(n5634), .Y(n4490) );
  CLKINVX1 U6309 ( .A(n5833), .Y(n4492) );
  CLKINVX1 U6310 ( .A(n5597), .Y(n4477) );
  NAND3X1 U6311 ( .A(n5998), .B(n6043), .C(n5876), .Y(n5467) );
  CLKINVX1 U6312 ( .A(n5392), .Y(n4513) );
  XNOR2X2 U6313 ( .A(n5991), .B(n6348), .Y(n5056) );
  NAND2X1 U6314 ( .A(n5469), .B(n5520), .Y(n5538) );
  XOR2X1 U6315 ( .A(n5061), .B(n5062), .Y(n5051) );
  XOR2X1 U6316 ( .A(n6349), .B(\add_0_root_add_0_root_add_92_2/carry[4] ), .Y(
        n5062) );
  NAND2X1 U6317 ( .A(n6004), .B(n4834), .Y(n4987) );
  NAND2X1 U6318 ( .A(n6350), .B(n4859), .Y(n5070) );
  NAND2X1 U6319 ( .A(n5153), .B(n6348), .Y(n4995) );
  CLKINVX1 U6320 ( .A(n5520), .Y(n4473) );
  NAND2X1 U6321 ( .A(n5991), .B(n4859), .Y(n5080) );
  NAND2BX1 U6322 ( .AN(n5089), .B(n5090), .Y(n5091) );
  NAND2BX1 U6323 ( .AN(n5092), .B(n5093), .Y(n5040) );
  NOR3X1 U6324 ( .A(n5053), .B(n5054), .C(n5055), .Y(n5052) );
  XOR2X1 U6325 ( .A(n5056), .B(n5057), .Y(n5055) );
  XOR2X1 U6326 ( .A(n5058), .B(n5059), .Y(n5053) );
  OA21XL U6327 ( .A0(n5092), .A1(n5926), .B0(n5093), .Y(n5924) );
  NAND2X1 U6328 ( .A(n6348), .B(n6350), .Y(n5926) );
  NAND3X1 U6329 ( .A(n6001), .B(n6053), .C(n5891), .Y(n5468) );
  NAND3X1 U6330 ( .A(n6060), .B(n6005), .C(n5553), .Y(n5469) );
  NAND2X1 U6331 ( .A(n6348), .B(n4834), .Y(n4973) );
  NAND2X1 U6332 ( .A(n5153), .B(n6004), .Y(n4992) );
  CLKINVX1 U6333 ( .A(n4911), .Y(n4847) );
  CLKINVX1 U6334 ( .A(n5079), .Y(n4542) );
  CLKINVX1 U6335 ( .A(n5076), .Y(n4548) );
  NOR2X1 U6336 ( .A(n6350), .B(n6348), .Y(n5041) );
  OA21XL U6337 ( .A0(n5041), .A1(n5092), .B0(n5093), .Y(n5088) );
  CLKINVX1 U6338 ( .A(n5016), .Y(n4469) );
  CLKBUFX3 U6339 ( .A(n6074), .Y(n6412) );
  CLKBUFX3 U6340 ( .A(n6074), .Y(n6413) );
  OAI31XL U6341 ( .A0(n5070), .A1(special_locate[2]), .A2(n4857), .B0(n4846), 
        .Y(n5069) );
  CLKINVX1 U6342 ( .A(isstring), .Y(n4845) );
  OAI2BB2XL U6343 ( .B0(n6298), .B1(n4986), .A0N(n6298), .A1N(pattern[55]), 
        .Y(n1390) );
  OAI2BB2XL U6344 ( .B0(n6298), .B1(n4983), .A0N(n6298), .A1N(pattern[52]), 
        .Y(n1393) );
  OAI2BB2XL U6345 ( .B0(n6298), .B1(n4985), .A0N(n6298), .A1N(pattern[54]), 
        .Y(n1391) );
  OAI2BB2XL U6346 ( .B0(n4456), .B1(n5033), .A0N(pattern_after[7]), .A1N(n4456), .Y(n1324) );
  OAI2BB2XL U6347 ( .B0(n4456), .B1(n5018), .A0N(pattern_after[0]), .A1N(n4456), .Y(n1373) );
  INVX3 U6348 ( .A(ispattern), .Y(n4846) );
  OAI32X4 U6349 ( .A0(n5011), .A1(n4649), .A2(n5012), .B0(n4449), .B1(n5013), 
        .Y(n4918) );
  AOI211X1 U6350 ( .A0(n4469), .A1(next_state[2]), .B0(n5014), .C0(n5015), .Y(
        n5013) );
  OAI21XL U6351 ( .A0(isstring), .A1(ispattern), .B0(n4849), .Y(n5047) );
  OAI211X1 U6352 ( .A0(n375), .A1(n4468), .B0(n6313), .C0(n4426), .Y(n5006) );
  NAND4X2 U6353 ( .A(n374), .B(n4993), .C(n4849), .D(n4468), .Y(n4989) );
  NOR4X1 U6354 ( .A(next_state[0]), .B(next_state[1]), .C(next_state[2]), .D(
        stringCounter[5]), .Y(n4948) );
  OAI221XL U6355 ( .A0(n5961), .A1(n4916), .B0(n6465), .B1(n5006), .C0(n5007), 
        .Y(n1379) );
  OAI221XL U6356 ( .A0(n5959), .A1(n4916), .B0(n6468), .B1(n5006), .C0(n5008), 
        .Y(n1377) );
  NOR2BX1 U6357 ( .AN(n4948), .B(stringCounter[4]), .Y(n4932) );
  NAND4X1 U6358 ( .A(n374), .B(n5977), .C(n4846), .D(n4849), .Y(n5042) );
  OAI2BB2XL U6359 ( .B0(n4464), .B1(n4986), .A0N(pattern[7]), .A1N(n4464), .Y(
        n1438) );
  OAI2BB2XL U6360 ( .B0(n4462), .B1(n4986), .A0N(n4462), .A1N(pattern[39]), 
        .Y(n1406) );
  OAI2BB2XL U6361 ( .B0(n4461), .B1(n4986), .A0N(n4461), .A1N(pattern[47]), 
        .Y(n1398) );
  OAI2BB2XL U6362 ( .B0(n4459), .B1(n4986), .A0N(n4459), .A1N(pattern[63]), 
        .Y(n1382) );
  OAI2BB2XL U6363 ( .B0(n4466), .B1(n4986), .A0N(n4466), .A1N(pattern[31]), 
        .Y(n1414) );
  OAI2BB2XL U6364 ( .B0(n4462), .B1(n4983), .A0N(n4462), .A1N(pattern[36]), 
        .Y(n1409) );
  OAI2BB2XL U6365 ( .B0(n4462), .B1(n4985), .A0N(n4462), .A1N(pattern[38]), 
        .Y(n1407) );
  OAI2BB2XL U6366 ( .B0(n4461), .B1(n4983), .A0N(n4461), .A1N(pattern[44]), 
        .Y(n1401) );
  OAI2BB2XL U6367 ( .B0(n4461), .B1(n4985), .A0N(n4461), .A1N(pattern[46]), 
        .Y(n1399) );
  OAI2BB2XL U6368 ( .B0(n4459), .B1(n4983), .A0N(n4459), .A1N(pattern[60]), 
        .Y(n1385) );
  OAI2BB2XL U6369 ( .B0(n4459), .B1(n4985), .A0N(n4459), .A1N(pattern[62]), 
        .Y(n1383) );
  OAI2BB2XL U6370 ( .B0(n4466), .B1(n4983), .A0N(n4466), .A1N(pattern[28]), 
        .Y(n1417) );
  OAI2BB2XL U6371 ( .B0(n4466), .B1(n4985), .A0N(n4466), .A1N(pattern[30]), 
        .Y(n1415) );
  OAI2BB2XL U6372 ( .B0(n4464), .B1(n4978), .A0N(pattern[0]), .A1N(n4464), .Y(
        n1445) );
  OAI2BB2XL U6373 ( .B0(n6300), .B1(n5027), .A0N(n5968), .A1N(n6300), .Y(n1364) );
  OAI2BB2XL U6374 ( .B0(n6300), .B1(n5031), .A0N(n5969), .A1N(n6300), .Y(n1336) );
  OAI2BB2XL U6375 ( .B0(n6300), .B1(n5029), .A0N(n5970), .A1N(n6300), .Y(n1350) );
  OAI2BB2XL U6376 ( .B0(n6300), .B1(n5028), .A0N(n5971), .A1N(n6300), .Y(n1358) );
  OAI222XL U6377 ( .A0(n5004), .A1(n6456), .B0(n6295), .B1(n5005), .C0(n5962), 
        .C1(n4916), .Y(n1381) );
  AOI2BB1X1 U6378 ( .A0N(n6350), .A1N(n6313), .B0(n4918), .Y(n5005) );
  OA21XL U6379 ( .A0(n6313), .A1(n5991), .B0(n5006), .Y(n5004) );
  AO22X1 U6380 ( .A0(chardata[5]), .A1(n4448), .B0(n6347), .B1(stringData[5]), 
        .Y(n1702) );
  OAI221XL U6381 ( .A0(n6349), .A1(n4915), .B0(n5960), .B1(n4916), .C0(n4917), 
        .Y(n1720) );
  AOI32XL U6382 ( .A0(n4918), .A1(n6349), .A2(\r720/carry[4] ), .B0(n4449), 
        .B1(n4919), .Y(n4917) );
  OA21XL U6383 ( .A0(n4426), .A1(\r720/carry[4] ), .B0(n4920), .Y(n4915) );
  OAI221X1 U6384 ( .A0(n6352), .A1(n4795), .B0(n6371), .B1(n4723), .C0(n5798), 
        .Y(n5583) );
  AOI22X1 U6385 ( .A0(n6358), .A1(stringData[112]), .B0(stringData[240]), .B1(
        n6365), .Y(n5798) );
  AOI22X1 U6386 ( .A0(n6359), .A1(stringData[116]), .B0(stringData[244]), .B1(
        n6364), .Y(n5754) );
  OAI221X1 U6387 ( .A0(n6352), .A1(n4789), .B0(n6277), .B1(n4717), .C0(n5809), 
        .Y(n5591) );
  AOI22X1 U6388 ( .A0(n6358), .A1(stringData[118]), .B0(stringData[246]), .B1(
        n6365), .Y(n5809) );
  OAI221X1 U6389 ( .A0(n6352), .A1(n4792), .B0(n6372), .B1(n4720), .C0(n5889), 
        .Y(n5816) );
  OAI221X1 U6390 ( .A0(n6352), .A1(n4794), .B0(n6371), .B1(n6009), .C0(n5881), 
        .Y(n5600) );
  AOI22X1 U6391 ( .A0(n6358), .A1(stringData[113]), .B0(stringData[241]), .B1(
        n6365), .Y(n5881) );
  OAI222X1 U6392 ( .A0(n5623), .A1(n6381), .B0(n5790), .B1(n6383), .C0(n6465), 
        .C1(n4636), .Y(n5720) );
  AOI221XL U6393 ( .A0(n6366), .A1(n4731), .B0(n6358), .B1(n4667), .C0(n5794), 
        .Y(n5790) );
  OAI22XL U6394 ( .A0(stringData[8]), .A1(n6370), .B0(stringData[136]), .B1(
        n6351), .Y(n5794) );
  OAI222X1 U6395 ( .A0(n5627), .A1(n6381), .B0(n5742), .B1(n6383), .C0(n6465), 
        .C1(n4643), .Y(n5696) );
  AOI221XL U6396 ( .A0(n6366), .A1(n4727), .B0(n6359), .B1(n4663), .C0(n5750), 
        .Y(n5742) );
  OAI22XL U6397 ( .A0(stringData[12]), .A1(n5655), .B0(stringData[140]), .B1(
        n6351), .Y(n5750) );
  AOI221XL U6398 ( .A0(n6366), .A1(n4724), .B0(n6359), .B1(n4660), .C0(n5761), 
        .Y(n5757) );
  OAI22XL U6399 ( .A0(stringData[15]), .A1(n6370), .B0(stringData[143]), .B1(
        n6351), .Y(n5761) );
  OAI222X1 U6400 ( .A0(n5615), .A1(n6381), .B0(n5801), .B1(n6383), .C0(n6465), 
        .C1(n4611), .Y(n5705) );
  AOI221XL U6401 ( .A0(n6366), .A1(n4725), .B0(n6359), .B1(n4661), .C0(n5805), 
        .Y(n5801) );
  OAI22XL U6402 ( .A0(stringData[14]), .A1(n5655), .B0(stringData[142]), .B1(
        n6351), .Y(n5805) );
  AOI221X1 U6403 ( .A0(n4743), .A1(n6355), .B0(n4679), .B1(n6375), .C0(n5751), 
        .Y(n5627) );
  OAI22XL U6404 ( .A0(stringData[108]), .A1(n6361), .B0(n6368), .B1(
        stringData[236]), .Y(n5751) );
  AOI221X1 U6405 ( .A0(n4744), .A1(n6355), .B0(n4680), .B1(n6377), .C0(n5887), 
        .Y(n5779) );
  OAI22XL U6406 ( .A0(stringData[107]), .A1(n6362), .B0(n6367), .B1(
        stringData[235]), .Y(n5887) );
  AOI221X1 U6407 ( .A0(n4741), .A1(n6355), .B0(n4677), .B1(n6378), .C0(n5806), 
        .Y(n5615) );
  OAI22XL U6408 ( .A0(stringData[110]), .A1(n6357), .B0(n6369), .B1(
        stringData[238]), .Y(n5806) );
  AOI221X1 U6409 ( .A0(n4746), .A1(n6355), .B0(n4682), .B1(n6377), .C0(n5883), 
        .Y(n5772) );
  OAI22XL U6410 ( .A0(stringData[105]), .A1(n6360), .B0(n6367), .B1(
        stringData[233]), .Y(n5883) );
  OAI222X1 U6411 ( .A0(n5772), .A1(n6381), .B0(n5773), .B1(n6383), .C0(n6465), 
        .C1(n4620), .Y(n5709) );
  AOI221XL U6412 ( .A0(n6366), .A1(n4730), .B0(n6358), .B1(n4666), .C0(n5774), 
        .Y(n5773) );
  OAI22XL U6413 ( .A0(stringData[9]), .A1(n5655), .B0(stringData[137]), .B1(
        n6351), .Y(n5774) );
  OAI222X1 U6414 ( .A0(n5779), .A1(n6381), .B0(n5780), .B1(n6383), .C0(n6465), 
        .C1(n4618), .Y(n5713) );
  AOI221XL U6415 ( .A0(n6366), .A1(n4728), .B0(n6358), .B1(n4664), .C0(n5781), 
        .Y(n5780) );
  OAI22XL U6416 ( .A0(stringData[11]), .A1(n5655), .B0(stringData[139]), .B1(
        n6351), .Y(n5781) );
  OAI221XL U6417 ( .A0(n6353), .A1(n4786), .B0(n6371), .B1(n5982), .C0(n5912), 
        .Y(n5860) );
  OAI221XL U6418 ( .A0(n6353), .A1(n4780), .B0(n6372), .B1(n4708), .C0(n5934), 
        .Y(n5759) );
  AOI22X1 U6419 ( .A0(n6358), .A1(stringData[127]), .B0(stringData[255]), .B1(
        n6365), .Y(n5934) );
  OAI221XL U6420 ( .A0(n6353), .A1(n4784), .B0(n6372), .B1(n4712), .C0(n5921), 
        .Y(n5852) );
  CLKINVX1 U6421 ( .A(n5763), .Y(n4638) );
  OAI221XL U6422 ( .A0(stringData[23]), .A1(n6304), .B0(n6473), .B1(n5587), 
        .C0(n5764), .Y(n5763) );
  AOI222XL U6423 ( .A0(n6305), .A1(n4804), .B0(n6306), .B1(n4772), .C0(n6307), 
        .C1(n4700), .Y(n5764) );
  CLKINVX1 U6424 ( .A(n5791), .Y(n4636) );
  OAI221XL U6425 ( .A0(stringData[24]), .A1(n6304), .B0(n6468), .B1(n5625), 
        .C0(n5792), .Y(n5791) );
  AOI222XL U6426 ( .A0(n6305), .A1(n4803), .B0(n6306), .B1(n4771), .C0(n6307), 
        .C1(n4699), .Y(n5792) );
  CLKINVX1 U6427 ( .A(n5859), .Y(n4620) );
  OAI221XL U6428 ( .A0(stringData[25]), .A1(n6304), .B0(n6473), .B1(n5860), 
        .C0(n5861), .Y(n5859) );
  AOI222XL U6429 ( .A0(n6305), .A1(n4802), .B0(n6306), .B1(n4770), .C0(n6307), 
        .C1(n4698), .Y(n5861) );
  CLKINVX1 U6430 ( .A(n5743), .Y(n4643) );
  OAI221XL U6431 ( .A0(stringData[28]), .A1(n6304), .B0(n6473), .B1(n5629), 
        .C0(n5745), .Y(n5743) );
  AOI222XL U6432 ( .A0(n6305), .A1(n4799), .B0(n6306), .B1(n4767), .C0(n6307), 
        .C1(n4695), .Y(n5745) );
  CLKINVX1 U6433 ( .A(n5802), .Y(n4611) );
  OAI221XL U6434 ( .A0(stringData[30]), .A1(n6304), .B0(n6468), .B1(n5803), 
        .C0(n5804), .Y(n5802) );
  CLKINVX1 U6435 ( .A(n5851), .Y(n4618) );
  OAI221XL U6436 ( .A0(stringData[27]), .A1(n6304), .B0(n6474), .B1(n5852), 
        .C0(n5853), .Y(n5851) );
  AOI222XL U6437 ( .A0(n6305), .A1(n4800), .B0(n6306), .B1(n4768), .C0(n6307), 
        .C1(n4696), .Y(n5853) );
  CLKINVX1 U6438 ( .A(n4995), .Y(n4832) );
  AOI211X1 U6439 ( .A0(n4829), .A1(n4552), .B0(n5101), .C0(n4518), .Y(n5100)
         );
  NOR3X2 U6440 ( .A(n4458), .B(reset), .C(n4911), .Y(n3297) );
  OAI32X1 U6441 ( .A0(n4846), .A1(patternCounter[2]), .A2(n4974), .B0(n4860), 
        .B1(n4975), .Y(n1447) );
  OAI32X1 U6442 ( .A0(n4846), .A1(n4976), .A2(n4974), .B0(n6021), .B1(n4977), 
        .Y(n1446) );
  OA21XL U6443 ( .A0(patternCounter[2]), .A1(n4846), .B0(n4975), .Y(n4977) );
  OAI32X1 U6444 ( .A0(n6004), .A1(ispattern), .A2(n4457), .B0(n6348), .B1(
        n4846), .Y(n1723) );
  XOR2X1 U6445 ( .A(n5424), .B(n4612), .Y(n5408) );
  XOR2X1 U6446 ( .A(n5357), .B(n5423), .Y(n5409) );
  OAI22XL U6447 ( .A0(pattern[0]), .A1(n4633), .B0(pattern[7]), .B1(n4615), 
        .Y(n5422) );
  OAI22XL U6448 ( .A0(stringCounter[0]), .A1(n4845), .B0(n4922), .B1(n4856), 
        .Y(n1717) );
  OAI22XL U6449 ( .A0(n6004), .A1(n4912), .B0(n6350), .B1(n4913), .Y(n1451) );
  OAI22XL U6450 ( .A0(n5960), .A1(n4449), .B0(n6349), .B1(n6313), .Y(n1721) );
  OAI22XL U6451 ( .A0(n5959), .A1(n4449), .B0(n6468), .B1(n6313), .Y(n1376) );
  OAI22XL U6452 ( .A0(n5958), .A1(n4449), .B0(n6476), .B1(n6313), .Y(n1374) );
  OAI22XL U6453 ( .A0(n5962), .A1(n4449), .B0(n6456), .B1(n6313), .Y(n1380) );
  OAI22XL U6454 ( .A0(n5961), .A1(n4449), .B0(n6464), .B1(n6313), .Y(n1378) );
  NAND4X1 U6455 ( .A(chardata[5]), .B(chardata[3]), .C(n5002), .D(n5003), .Y(
        n4971) );
  NOR4X1 U6456 ( .A(chardata[7]), .B(chardata[6]), .C(chardata[4]), .D(
        chardata[2]), .Y(n5003) );
  NOR2X1 U6457 ( .A(chardata[0]), .B(n6393), .Y(n5002) );
  AOI22X1 U6458 ( .A0(n6359), .A1(stringData[120]), .B0(stringData[248]), .B1(
        n6364), .Y(n5793) );
  NAND4X1 U6459 ( .A(n4829), .B(n5154), .C(patternCounter[3]), .D(n4860), .Y(
        n5139) );
  OAI31XL U6460 ( .A0(n5155), .A1(n5131), .A2(n5102), .B0(n5156), .Y(n5154) );
  NAND4X1 U6461 ( .A(n5157), .B(n5158), .C(n5159), .D(n5160), .Y(n5156) );
  XOR2X1 U6462 ( .A(n5262), .B(n5108), .Y(n5157) );
  OAI2BB2XL U6463 ( .B0(n4853), .B1(n4922), .A0N(N1245), .A1N(isstring), .Y(
        n1711) );
  OAI2BB2XL U6464 ( .B0(n4854), .B1(n4922), .A0N(N1244), .A1N(isstring), .Y(
        n1713) );
  OAI2BB2XL U6465 ( .B0(n4855), .B1(n4922), .A0N(N1243), .A1N(isstring), .Y(
        n1715) );
  OAI2BB2XL U6466 ( .B0(n4851), .B1(n4922), .A0N(N1246), .A1N(isstring), .Y(
        n1709) );
  OAI221X1 U6467 ( .A0(n6352), .A1(n4788), .B0(n6372), .B1(n4716), .C0(n5765), 
        .Y(n5587) );
  AOI2BB2X1 U6468 ( .B0(stringData[247]), .B1(n6365), .A0N(n6362), .A1N(n6007), 
        .Y(n5765) );
  CLKINVX1 U6469 ( .A(n5758), .Y(n4616) );
  OAI221XL U6470 ( .A0(stringData[31]), .A1(n6304), .B0(n6473), .B1(n5759), 
        .C0(n5760), .Y(n5758) );
  AOI222XL U6471 ( .A0(n6305), .A1(n4796), .B0(n6306), .B1(n4764), .C0(n6307), 
        .C1(n4692), .Y(n5760) );
  CLKINVX1 U6472 ( .A(n5796), .Y(n4635) );
  OAI221XL U6473 ( .A0(stringData[16]), .A1(n6304), .B0(n6473), .B1(n5583), 
        .C0(n5797), .Y(n5796) );
  AOI222XL U6474 ( .A0(n6305), .A1(n4811), .B0(n6306), .B1(n4779), .C0(n6307), 
        .C1(n4707), .Y(n5797) );
  CLKINVX1 U6475 ( .A(n5776), .Y(n4625) );
  OAI221XL U6476 ( .A0(stringData[17]), .A1(n6304), .B0(n6468), .B1(n5600), 
        .C0(n5777), .Y(n5776) );
  AOI222XL U6477 ( .A0(n6305), .A1(n4810), .B0(n6306), .B1(n4778), .C0(n6307), 
        .C1(n4706), .Y(n5777) );
  OAI221XL U6478 ( .A0(stringData[20]), .A1(n6304), .B0(n6473), .B1(n5575), 
        .C0(n5753), .Y(n5752) );
  AOI222XL U6479 ( .A0(n6305), .A1(n4807), .B0(n6306), .B1(n4775), .C0(n6307), 
        .C1(n4703), .Y(n5753) );
  CLKINVX1 U6480 ( .A(n5815), .Y(n4624) );
  OAI221XL U6481 ( .A0(stringData[19]), .A1(n6304), .B0(n6474), .B1(n5816), 
        .C0(n5817), .Y(n5815) );
  AOI222XL U6482 ( .A0(n6305), .A1(n4808), .B0(n6306), .B1(n4776), .C0(n6307), 
        .C1(n4704), .Y(n5817) );
  OAI221XL U6483 ( .A0(stringData[22]), .A1(n6304), .B0(n6468), .B1(n5591), 
        .C0(n5808), .Y(n5807) );
  AOI222XL U6484 ( .A0(n6305), .A1(n4805), .B0(n6306), .B1(n4773), .C0(n6307), 
        .C1(n4701), .Y(n5808) );
  OAI2BB2XL U6485 ( .B0(n6393), .B1(n6317), .A0N(n6317), .A1N(stringData[241]), 
        .Y(n1466) );
  OAI2BB2XL U6486 ( .B0(n6393), .B1(n6316), .A0N(n6316), .A1N(stringData[249]), 
        .Y(n1458) );
  OAI2BB2XL U6487 ( .B0(n6393), .B1(n6330), .A0N(n6330), .A1N(stringData[137]), 
        .Y(n1570) );
  OAI2BB2XL U6488 ( .B0(n6393), .B1(n6345), .A0N(n6345), .A1N(stringData[17]), 
        .Y(n1690) );
  OAI2BB2XL U6489 ( .B0(n6393), .B1(n6344), .A0N(n6344), .A1N(stringData[25]), 
        .Y(n1682) );
  OAI2BB2XL U6490 ( .B0(n6393), .B1(n6333), .A0N(n6333), .A1N(stringData[113]), 
        .Y(n1594) );
  OAI2BB2XL U6491 ( .B0(n6393), .B1(n6332), .A0N(n6332), .A1N(stringData[121]), 
        .Y(n1586) );
  OAI2BB2XL U6492 ( .B0(n6393), .B1(n6346), .A0N(n6346), .A1N(stringData[9]), 
        .Y(n1698) );
  OAI2BB2XL U6493 ( .B0(n6393), .B1(n6343), .A0N(n6343), .A1N(stringData[33]), 
        .Y(n1674) );
  OAI2BB2XL U6494 ( .B0(n6393), .B1(n6335), .A0N(n6335), .A1N(stringData[97]), 
        .Y(n1610) );
  OAI2BB2XL U6495 ( .B0(n6391), .B1(n6317), .A0N(n6317), .A1N(stringData[240]), 
        .Y(n1467) );
  OAI2BB2XL U6496 ( .B0(n6395), .B1(n6317), .A0N(n6317), .A1N(stringData[242]), 
        .Y(n1465) );
  OAI2BB2XL U6497 ( .B0(n6397), .B1(n6317), .A0N(n6317), .A1N(stringData[243]), 
        .Y(n1464) );
  OAI2BB2XL U6498 ( .B0(n6399), .B1(n6317), .A0N(n6317), .A1N(stringData[244]), 
        .Y(n1463) );
  OAI2BB2XL U6499 ( .B0(n6401), .B1(n6317), .A0N(n6317), .A1N(stringData[245]), 
        .Y(n1462) );
  OAI2BB2XL U6500 ( .B0(n6403), .B1(n6317), .A0N(n6317), .A1N(stringData[246]), 
        .Y(n1461) );
  OAI2BB2XL U6501 ( .B0(n6405), .B1(n6317), .A0N(n6317), .A1N(stringData[247]), 
        .Y(n1460) );
  OAI2BB2XL U6502 ( .B0(n6391), .B1(n6316), .A0N(n6316), .A1N(stringData[248]), 
        .Y(n1459) );
  OAI2BB2XL U6503 ( .B0(n6395), .B1(n6316), .A0N(n6316), .A1N(stringData[250]), 
        .Y(n1457) );
  OAI2BB2XL U6504 ( .B0(n6397), .B1(n6316), .A0N(n6316), .A1N(stringData[251]), 
        .Y(n1456) );
  OAI2BB2XL U6505 ( .B0(n6399), .B1(n6316), .A0N(n6316), .A1N(stringData[252]), 
        .Y(n1455) );
  OAI2BB2XL U6506 ( .B0(n6401), .B1(n6316), .A0N(n6316), .A1N(stringData[253]), 
        .Y(n1454) );
  OAI2BB2XL U6507 ( .B0(n6403), .B1(n6316), .A0N(n6316), .A1N(stringData[254]), 
        .Y(n1453) );
  OAI2BB2XL U6508 ( .B0(n6405), .B1(n6316), .A0N(n6316), .A1N(stringData[255]), 
        .Y(n1452) );
  OAI2BB2XL U6509 ( .B0(n6391), .B1(n6330), .A0N(n6330), .A1N(stringData[136]), 
        .Y(n1571) );
  OAI2BB2XL U6510 ( .B0(n6395), .B1(n6330), .A0N(n6330), .A1N(stringData[138]), 
        .Y(n1569) );
  OAI2BB2XL U6511 ( .B0(n6397), .B1(n6330), .A0N(n6330), .A1N(stringData[139]), 
        .Y(n1568) );
  OAI2BB2XL U6512 ( .B0(n6399), .B1(n6330), .A0N(n6330), .A1N(stringData[140]), 
        .Y(n1567) );
  OAI2BB2XL U6513 ( .B0(n6401), .B1(n6330), .A0N(n6330), .A1N(stringData[141]), 
        .Y(n1566) );
  OAI2BB2XL U6514 ( .B0(n6403), .B1(n6330), .A0N(n6330), .A1N(stringData[142]), 
        .Y(n1565) );
  OAI2BB2XL U6515 ( .B0(n6405), .B1(n6330), .A0N(n6330), .A1N(stringData[143]), 
        .Y(n1564) );
  OAI2BB2XL U6516 ( .B0(n6391), .B1(n6345), .A0N(n6345), .A1N(stringData[16]), 
        .Y(n1691) );
  OAI2BB2XL U6517 ( .B0(n6395), .B1(n6345), .A0N(n6345), .A1N(stringData[18]), 
        .Y(n1689) );
  OAI2BB2XL U6518 ( .B0(n6397), .B1(n6345), .A0N(n6345), .A1N(stringData[19]), 
        .Y(n1688) );
  OAI2BB2XL U6519 ( .B0(n6399), .B1(n6345), .A0N(n6345), .A1N(stringData[20]), 
        .Y(n1687) );
  OAI2BB2XL U6520 ( .B0(n6401), .B1(n6345), .A0N(n6345), .A1N(stringData[21]), 
        .Y(n1686) );
  OAI2BB2XL U6521 ( .B0(n6403), .B1(n6345), .A0N(n6345), .A1N(stringData[22]), 
        .Y(n1685) );
  OAI2BB2XL U6522 ( .B0(n6405), .B1(n6345), .A0N(n6345), .A1N(stringData[23]), 
        .Y(n1684) );
  OAI2BB2XL U6523 ( .B0(n6391), .B1(n6344), .A0N(n6344), .A1N(stringData[24]), 
        .Y(n1683) );
  OAI2BB2XL U6524 ( .B0(n6395), .B1(n6344), .A0N(n6344), .A1N(stringData[26]), 
        .Y(n1681) );
  OAI2BB2XL U6525 ( .B0(n6397), .B1(n6344), .A0N(n6344), .A1N(stringData[27]), 
        .Y(n1680) );
  OAI2BB2XL U6526 ( .B0(n6399), .B1(n6344), .A0N(n6344), .A1N(stringData[28]), 
        .Y(n1679) );
  OAI2BB2XL U6527 ( .B0(n6401), .B1(n6344), .A0N(n6344), .A1N(stringData[29]), 
        .Y(n1678) );
  OAI2BB2XL U6528 ( .B0(n6403), .B1(n6344), .A0N(n6344), .A1N(stringData[30]), 
        .Y(n1677) );
  OAI2BB2XL U6529 ( .B0(n6405), .B1(n6344), .A0N(n6344), .A1N(stringData[31]), 
        .Y(n1676) );
  OAI2BB2XL U6530 ( .B0(n6391), .B1(n6333), .A0N(n6333), .A1N(stringData[112]), 
        .Y(n1595) );
  OAI2BB2XL U6531 ( .B0(n6395), .B1(n6333), .A0N(n6333), .A1N(stringData[114]), 
        .Y(n1593) );
  OAI2BB2XL U6532 ( .B0(n6397), .B1(n6333), .A0N(n6333), .A1N(stringData[115]), 
        .Y(n1592) );
  OAI2BB2XL U6533 ( .B0(n6399), .B1(n6333), .A0N(n6333), .A1N(stringData[116]), 
        .Y(n1591) );
  OAI2BB2XL U6534 ( .B0(n6401), .B1(n6333), .A0N(n6333), .A1N(stringData[117]), 
        .Y(n1590) );
  OAI2BB2XL U6535 ( .B0(n6403), .B1(n6333), .A0N(n6333), .A1N(stringData[118]), 
        .Y(n1589) );
  OAI2BB2XL U6536 ( .B0(n6405), .B1(n6333), .A0N(n6333), .A1N(stringData[119]), 
        .Y(n1588) );
  OAI2BB2XL U6537 ( .B0(n6391), .B1(n6332), .A0N(n6332), .A1N(stringData[120]), 
        .Y(n1587) );
  OAI2BB2XL U6538 ( .B0(n6395), .B1(n6332), .A0N(n6332), .A1N(stringData[122]), 
        .Y(n1585) );
  OAI2BB2XL U6539 ( .B0(n6397), .B1(n6332), .A0N(n6332), .A1N(stringData[123]), 
        .Y(n1584) );
  OAI2BB2XL U6540 ( .B0(n6399), .B1(n6332), .A0N(n6332), .A1N(stringData[124]), 
        .Y(n1583) );
  OAI2BB2XL U6541 ( .B0(n6401), .B1(n6332), .A0N(n6332), .A1N(stringData[125]), 
        .Y(n1582) );
  OAI2BB2XL U6542 ( .B0(n6403), .B1(n6332), .A0N(n6332), .A1N(stringData[126]), 
        .Y(n1581) );
  OAI2BB2XL U6543 ( .B0(n6405), .B1(n6332), .A0N(n6332), .A1N(stringData[127]), 
        .Y(n1580) );
  OAI2BB2XL U6544 ( .B0(n6391), .B1(n6346), .A0N(n6346), .A1N(stringData[8]), 
        .Y(n1699) );
  OAI2BB2XL U6545 ( .B0(n6395), .B1(n6346), .A0N(n6346), .A1N(stringData[10]), 
        .Y(n1697) );
  OAI2BB2XL U6546 ( .B0(n6397), .B1(n6346), .A0N(n6346), .A1N(stringData[11]), 
        .Y(n1696) );
  OAI2BB2XL U6547 ( .B0(n6399), .B1(n6346), .A0N(n6346), .A1N(stringData[12]), 
        .Y(n1695) );
  OAI2BB2XL U6548 ( .B0(n6401), .B1(n6346), .A0N(n6346), .A1N(stringData[13]), 
        .Y(n1694) );
  OAI2BB2XL U6549 ( .B0(n6403), .B1(n6346), .A0N(n6346), .A1N(stringData[14]), 
        .Y(n1693) );
  OAI2BB2XL U6550 ( .B0(n6405), .B1(n6346), .A0N(n6346), .A1N(stringData[15]), 
        .Y(n1692) );
  OAI2BB2XL U6551 ( .B0(n6391), .B1(n6343), .A0N(n6343), .A1N(stringData[32]), 
        .Y(n1675) );
  OAI2BB2XL U6552 ( .B0(n6395), .B1(n6343), .A0N(n6343), .A1N(stringData[34]), 
        .Y(n1673) );
  OAI2BB2XL U6553 ( .B0(n6397), .B1(n6343), .A0N(n6343), .A1N(stringData[35]), 
        .Y(n1672) );
  OAI2BB2XL U6554 ( .B0(n6399), .B1(n6343), .A0N(n6343), .A1N(stringData[36]), 
        .Y(n1671) );
  OAI2BB2XL U6555 ( .B0(n6401), .B1(n6343), .A0N(n6343), .A1N(stringData[37]), 
        .Y(n1670) );
  OAI2BB2XL U6556 ( .B0(n6403), .B1(n6343), .A0N(n6343), .A1N(stringData[38]), 
        .Y(n1669) );
  OAI2BB2XL U6557 ( .B0(n6405), .B1(n6343), .A0N(n6343), .A1N(stringData[39]), 
        .Y(n1668) );
  OAI2BB2XL U6558 ( .B0(n6391), .B1(n6335), .A0N(n6335), .A1N(stringData[96]), 
        .Y(n1611) );
  OAI2BB2XL U6559 ( .B0(n6395), .B1(n6335), .A0N(n6335), .A1N(stringData[98]), 
        .Y(n1609) );
  OAI2BB2XL U6560 ( .B0(n6397), .B1(n6335), .A0N(n6335), .A1N(stringData[99]), 
        .Y(n1608) );
  OAI2BB2XL U6561 ( .B0(n6399), .B1(n6335), .A0N(n6335), .A1N(stringData[100]), 
        .Y(n1607) );
  OAI2BB2XL U6562 ( .B0(n6401), .B1(n6335), .A0N(n6335), .A1N(stringData[101]), 
        .Y(n1606) );
  OAI2BB2XL U6563 ( .B0(n6403), .B1(n6335), .A0N(n6335), .A1N(stringData[102]), 
        .Y(n1605) );
  OAI2BB2XL U6564 ( .B0(n6405), .B1(n6335), .A0N(n6335), .A1N(stringData[103]), 
        .Y(n1604) );
  OA21XL U6565 ( .A0(patternCounter[1]), .A1(n4846), .B0(n4972), .Y(n4975) );
  OAI32X1 U6566 ( .A0(n4845), .A1(stringCounter[5]), .A2(n4852), .B0(n4921), 
        .B1(n4850), .Y(n1719) );
  CLKINVX1 U6567 ( .A(\add_802_S2/carry[5] ), .Y(n4852) );
  OA21XL U6568 ( .A0(\add_802_S2/carry[5] ), .A1(n4845), .B0(n4922), .Y(n4921)
         );
  OAI221X1 U6569 ( .A0(n6352), .A1(n4790), .B0(n6371), .B1(n4718), .C0(n5903), 
        .Y(n5822) );
  OAI221X1 U6570 ( .A0(n6352), .A1(n4793), .B0(n6371), .B1(n4721), .C0(n5895), 
        .Y(n5830) );
  AOI221X1 U6571 ( .A0(n4747), .A1(n6355), .B0(n4683), .B1(n6375), .C0(n5795), 
        .Y(n5623) );
  OAI22XL U6572 ( .A0(stringData[104]), .A1(n6361), .B0(n6369), .B1(
        stringData[232]), .Y(n5795) );
  AOI221X1 U6573 ( .A0(n4740), .A1(n6355), .B0(n4676), .B1(n6377), .C0(n5762), 
        .Y(n5619) );
  OAI22XL U6574 ( .A0(stringData[111]), .A1(n6361), .B0(n6369), .B1(
        stringData[239]), .Y(n5762) );
  AOI221X1 U6575 ( .A0(n4742), .A1(n6356), .B0(n4678), .B1(n6377), .C0(n5900), 
        .Y(n5783) );
  OAI22XL U6576 ( .A0(stringData[109]), .A1(n6360), .B0(n6368), .B1(
        stringData[237]), .Y(n5900) );
  AOI221X1 U6577 ( .A0(n4745), .A1(n6355), .B0(n4681), .B1(n6377), .C0(n5893), 
        .Y(n5787) );
  OAI22XL U6578 ( .A0(stringData[106]), .A1(n6360), .B0(n6369), .B1(
        stringData[234]), .Y(n5893) );
  AOI211X1 U6579 ( .A0(n4660), .A1(n6378), .B0(n6366), .C0(n5935), .Y(n5620)
         );
  OAI22XL U6580 ( .A0(stringData[207]), .A1(n6349), .B0(stringData[143]), .B1(
        n6476), .Y(n5935) );
  AOI211X1 U6581 ( .A0(n4661), .A1(n6378), .B0(n6366), .C0(n5957), .Y(n5616)
         );
  OAI22XL U6582 ( .A0(stringData[206]), .A1(n6349), .B0(stringData[142]), .B1(
        n6476), .Y(n5957) );
  AOI211X1 U6583 ( .A0(n4662), .A1(n6375), .B0(n6366), .C0(n5899), .Y(n5545)
         );
  OAI22XL U6584 ( .A0(stringData[205]), .A1(n6349), .B0(stringData[141]), .B1(
        n6476), .Y(n5899) );
  AOI211X1 U6585 ( .A0(n4666), .A1(n6378), .B0(n6366), .C0(n5913), .Y(n5858)
         );
  OAI22XL U6586 ( .A0(stringData[201]), .A1(n6349), .B0(stringData[137]), .B1(
        n6477), .Y(n5913) );
  AOI211X1 U6587 ( .A0(n4665), .A1(n6376), .B0(n6366), .C0(n5947), .Y(n5844)
         );
  OAI22XL U6588 ( .A0(stringData[202]), .A1(n6349), .B0(stringData[138]), .B1(
        n6476), .Y(n5947) );
  OAI222X1 U6589 ( .A0(n5787), .A1(n6381), .B0(n5788), .B1(n6383), .C0(n6465), 
        .C1(n4613), .Y(n5733) );
  AOI221XL U6590 ( .A0(n6366), .A1(n4729), .B0(n6359), .B1(n4665), .C0(n5789), 
        .Y(n5788) );
  OAI22XL U6591 ( .A0(stringData[10]), .A1(n5655), .B0(stringData[138]), .B1(
        n6351), .Y(n5789) );
  OAI221XL U6592 ( .A0(n6353), .A1(n4785), .B0(n6372), .B1(n4713), .C0(n5946), 
        .Y(n5846) );
  OAI221XL U6593 ( .A0(n6352), .A1(n4782), .B0(n6371), .B1(n4710), .C0(n5898), 
        .Y(n5835) );
  OAI222X1 U6594 ( .A0(n5783), .A1(n6381), .B0(n5784), .B1(n6383), .C0(n6465), 
        .C1(n4622), .Y(n5725) );
  AOI221XL U6595 ( .A0(n6366), .A1(n4726), .B0(n6358), .B1(n4662), .C0(n5785), 
        .Y(n5784) );
  OAI22XL U6596 ( .A0(stringData[13]), .A1(n5655), .B0(stringData[141]), .B1(
        n6351), .Y(n5785) );
  OAI222XL U6597 ( .A0(n4629), .A1(n6381), .B0(n5727), .B1(n6383), .C0(n6465), 
        .C1(n4621), .Y(n5726) );
  AOI221XL U6598 ( .A0(n6366), .A1(n4734), .B0(n6359), .B1(n4670), .C0(n5728), 
        .Y(n5727) );
  OAI22XL U6599 ( .A0(stringData[5]), .A1(n5655), .B0(stringData[133]), .B1(
        n6351), .Y(n5728) );
  OA21XL U6600 ( .A0(n5373), .A1(n5981), .B0(n5736), .Y(n5683) );
  AOI221XL U6601 ( .A0(pattern_after[12]), .A1(n4639), .B0(pattern_after[15]), 
        .B1(n4614), .C0(n5447), .Y(n5684) );
  OAI32X1 U6602 ( .A0(n5737), .A1(n5738), .A2(n5739), .B0(n5740), .B1(n5741), 
        .Y(n5736) );
  XOR2X1 U6603 ( .A(n5875), .B(n5202), .Y(n5603) );
  XOR2X1 U6604 ( .A(n5869), .B(n5204), .Y(n5604) );
  AOI221XL U6605 ( .A0(pattern_after[36]), .A1(n4569), .B0(n5974), .B1(n4563), 
        .C0(n5607), .Y(n5606) );
  NAND4X1 U6606 ( .A(n5663), .B(n5664), .C(n5665), .D(n5666), .Y(n5445) );
  XOR2X1 U6607 ( .A(n5824), .B(n4594), .Y(n5663) );
  XOR2X1 U6608 ( .A(n5818), .B(n4577), .Y(n5664) );
  AOI221XL U6609 ( .A0(pattern_after[20]), .A1(n4567), .B0(pattern_after[22]), 
        .B1(n4597), .C0(n5667), .Y(n5666) );
  XOR2X1 U6610 ( .A(n5848), .B(n4584), .Y(n5638) );
  XOR2X1 U6611 ( .A(n5854), .B(n5221), .Y(n5637) );
  AOI221XL U6612 ( .A0(pattern_after[28]), .A1(n4568), .B0(n5975), .B1(n4562), 
        .C0(n5641), .Y(n5640) );
  OAI22XL U6613 ( .A0(patternCounter[1]), .A1(n5086), .B0(n6348), .B1(n5084), 
        .Y(n5101) );
  OAI22XL U6614 ( .A0(pattern_after[0]), .A1(n4633), .B0(pattern_after[7]), 
        .B1(n4615), .Y(n5716) );
  NAND4X1 U6615 ( .A(n5563), .B(n5564), .C(n5565), .D(n5566), .Y(n5443) );
  XOR2X1 U6616 ( .A(n5890), .B(n5187), .Y(n5564) );
  XOR2X1 U6617 ( .A(n5896), .B(n4573), .Y(n5563) );
  AOI221XL U6618 ( .A0(pattern_after[46]), .A1(n4600), .B0(pattern_after[47]), 
        .B1(n4590), .C0(n5567), .Y(n5566) );
  NAND4X1 U6619 ( .A(n5685), .B(n5686), .C(n5687), .D(n5688), .Y(n5447) );
  AOI222XL U6620 ( .A0(pattern_after[0]), .A1(n4633), .B0(n5716), .B1(n5695), 
        .C0(pattern_after[7]), .C1(n4615), .Y(n5687) );
  CLKINVX1 U6621 ( .A(n5799), .Y(n4634) );
  OAI221XL U6622 ( .A0(stringData[160]), .A1(n6352), .B0(stringData[32]), .B1(
        n6277), .C0(n5800), .Y(n5799) );
  AOI2BB2X1 U6623 ( .B0(n6364), .B1(n4827), .A0N(stringData[96]), .A1N(n6362), 
        .Y(n5800) );
  CLKINVX1 U6624 ( .A(n5755), .Y(n4641) );
  OAI221XL U6625 ( .A0(stringData[164]), .A1(n6351), .B0(stringData[36]), .B1(
        n5655), .C0(n5756), .Y(n5755) );
  AOI2BB2X1 U6626 ( .B0(n6364), .B1(n4823), .A0N(stringData[100]), .A1N(n6362), 
        .Y(n5756) );
  CLKINVX1 U6627 ( .A(n5873), .Y(n4627) );
  OAI221XL U6628 ( .A0(stringData[163]), .A1(n6351), .B0(stringData[35]), .B1(
        n6371), .C0(n5874), .Y(n5873) );
  AOI2BB2X1 U6629 ( .B0(n6364), .B1(n4824), .A0N(stringData[99]), .A1N(n6362), 
        .Y(n5874) );
  CLKINVX1 U6630 ( .A(n5810), .Y(n4630) );
  OAI221XL U6631 ( .A0(stringData[166]), .A1(n6352), .B0(stringData[38]), .B1(
        n5655), .C0(n5811), .Y(n5810) );
  AOI2BB2X1 U6632 ( .B0(n6364), .B1(n4821), .A0N(stringData[102]), .A1N(n6362), 
        .Y(n5811) );
  CLKINVX1 U6633 ( .A(n5879), .Y(n4626) );
  OAI221XL U6634 ( .A0(stringData[161]), .A1(n6351), .B0(stringData[33]), .B1(
        n6371), .C0(n5880), .Y(n5879) );
  AOI2BB2X1 U6635 ( .B0(n6364), .B1(n4826), .A0N(stringData[97]), .A1N(n6362), 
        .Y(n5880) );
  CLKINVX1 U6636 ( .A(n5867), .Y(n4628) );
  OAI221XL U6637 ( .A0(stringData[162]), .A1(n6351), .B0(stringData[34]), .B1(
        n6371), .C0(n5868), .Y(n5867) );
  AOI2BB2X1 U6638 ( .B0(n6364), .B1(n4825), .A0N(stringData[98]), .A1N(n6362), 
        .Y(n5868) );
  CLKINVX1 U6639 ( .A(n5838), .Y(n4629) );
  OAI221XL U6640 ( .A0(stringData[165]), .A1(n6352), .B0(stringData[37]), .B1(
        n5655), .C0(n5839), .Y(n5838) );
  AOI2BB2X1 U6641 ( .B0(n6364), .B1(n4822), .A0N(stringData[101]), .A1N(n6362), 
        .Y(n5839) );
  CLKINVX1 U6642 ( .A(n5766), .Y(n4637) );
  OAI221XL U6643 ( .A0(stringData[167]), .A1(n6351), .B0(stringData[39]), .B1(
        n6277), .C0(n5767), .Y(n5766) );
  AOI2BB2X1 U6644 ( .B0(n6364), .B1(n4820), .A0N(stringData[103]), .A1N(n6362), 
        .Y(n5767) );
  CLKINVX1 U6645 ( .A(n5821), .Y(n4621) );
  OAI221XL U6646 ( .A0(stringData[21]), .A1(n6304), .B0(n6474), .B1(n5822), 
        .C0(n5823), .Y(n5821) );
  AOI222XL U6647 ( .A0(n6305), .A1(n4806), .B0(n6306), .B1(n4774), .C0(n6307), 
        .C1(n4702), .Y(n5823) );
  CLKINVX1 U6648 ( .A(n5845), .Y(n4613) );
  OAI221XL U6649 ( .A0(stringData[26]), .A1(n6304), .B0(n6474), .B1(n5846), 
        .C0(n5847), .Y(n5845) );
  AOI222XL U6650 ( .A0(n6305), .A1(n4801), .B0(n6306), .B1(n4769), .C0(n6307), 
        .C1(n4697), .Y(n5847) );
  CLKINVX1 U6651 ( .A(n5834), .Y(n4622) );
  OAI221XL U6652 ( .A0(stringData[29]), .A1(n6304), .B0(n6474), .B1(n5835), 
        .C0(n5836), .Y(n5834) );
  AOI222XL U6653 ( .A0(n6305), .A1(n4798), .B0(n6306), .B1(n4766), .C0(n6307), 
        .C1(n4694), .Y(n5836) );
  CLKINVX1 U6654 ( .A(n5829), .Y(n4623) );
  OAI221XL U6655 ( .A0(stringData[18]), .A1(n6304), .B0(n6474), .B1(n5830), 
        .C0(n5831), .Y(n5829) );
  AOI222XL U6656 ( .A0(n6305), .A1(n4809), .B0(n6306), .B1(n4777), .C0(n6307), 
        .C1(n4705), .Y(n5831) );
  CLKBUFX3 U6657 ( .A(n6479), .Y(n6451) );
  AND2X2 U6658 ( .A(n5514), .B(n5515), .Y(n5440) );
  AOI211X1 U6659 ( .A0(pattern_after[54]), .A1(n4596), .B0(n5516), .C0(n5517), 
        .Y(n5515) );
  NOR4X1 U6660 ( .A(n5533), .B(n5534), .C(n5535), .D(n5536), .Y(n5514) );
  OAI32X1 U6661 ( .A0(n4596), .A1(pattern_after[54]), .A2(n4473), .B0(n5518), 
        .B1(n6067), .Y(n5517) );
  OAI211X1 U6662 ( .A0(stringData[85]), .A1(n6372), .B0(n6369), .C0(n5902), 
        .Y(n5513) );
  OAI211X1 U6663 ( .A0(stringData[81]), .A1(n6372), .B0(n6369), .C0(n5907), 
        .Y(n5602) );
  OAI211X1 U6664 ( .A0(stringData[84]), .A1(n6372), .B0(n6369), .C0(n5660), 
        .Y(n5508) );
  OAI211X1 U6665 ( .A0(stringData[80]), .A1(n6372), .B0(n6369), .C0(n5657), 
        .Y(n5503) );
  OAI211X1 U6666 ( .A0(stringData[86]), .A1(n6372), .B0(n6369), .C0(n5951), 
        .Y(n5593) );
  OAI211X1 U6667 ( .A0(stringData[82]), .A1(n6372), .B0(n6369), .C0(n5941), 
        .Y(n5866) );
  OAI211X1 U6668 ( .A0(stringData[83]), .A1(n6372), .B0(n6369), .C0(n5916), 
        .Y(n5872) );
  AOI2BB2X1 U6669 ( .B0(n4776), .B1(match_index[4]), .A0N(stringData[147]), 
        .A1N(n6476), .Y(n5916) );
  AOI211X1 U6670 ( .A0(n4700), .A1(n6376), .B0(n6366), .C0(n5937), .Y(n5588)
         );
  OAI22XL U6671 ( .A0(stringData[215]), .A1(n6349), .B0(stringData[151]), .B1(
        n6476), .Y(n5937) );
  AOI211X1 U6672 ( .A0(n4667), .A1(n6378), .B0(n6366), .C0(n5671), .Y(n5561)
         );
  OAI22XL U6673 ( .A0(stringData[200]), .A1(n6349), .B0(stringData[136]), .B1(
        n6477), .Y(n5671) );
  AOI211X1 U6674 ( .A0(n4664), .A1(n6378), .B0(n6366), .C0(n5922), .Y(n5850)
         );
  OAI22XL U6675 ( .A0(stringData[203]), .A1(n6349), .B0(stringData[139]), .B1(
        n6476), .Y(n5922) );
  AOI211X1 U6676 ( .A0(n4663), .A1(n6376), .B0(n6366), .C0(n5675), .Y(n5529)
         );
  OAI22XL U6677 ( .A0(stringData[204]), .A1(n6349), .B0(stringData[140]), .B1(
        n6477), .Y(n5675) );
  NAND4X2 U6678 ( .A(pattern[5]), .B(n5425), .C(n6010), .D(n5983), .Y(n5417)
         );
  AOI22X1 U6679 ( .A0(stringData[101]), .A1(n6303), .B0(n5820), .B1(n6468), 
        .Y(n5901) );
  OAI222XL U6680 ( .A0(n5642), .A1(n6045), .B0(n4492), .B1(n5643), .C0(n5644), 
        .C1(n6000), .Y(n5641) );
  AOI221XL U6681 ( .A0(n5645), .A1(n6038), .B0(n5248), .B1(n5993), .C0(n5646), 
        .Y(n5643) );
  OAI22XL U6682 ( .A0(pattern_after[31]), .A1(n4588), .B0(pattern_after[30]), 
        .B1(n4598), .Y(n5646) );
  NAND4X1 U6683 ( .A(pattern[6]), .B(pattern[4]), .C(n5425), .D(n6008), .Y(
        n5012) );
  AOI2BB1X1 U6684 ( .A0N(n4562), .A1N(n5309), .B0(pattern[24]), .Y(n5243) );
  OAI22XL U6685 ( .A0(pattern_after[15]), .A1(n4614), .B0(pattern_after[12]), 
        .B1(n4639), .Y(n5739) );
  OAI22XL U6686 ( .A0(pattern_after[14]), .A1(n4608), .B0(pattern_after[8]), 
        .B1(n4632), .Y(n5738) );
  OAI222XL U6687 ( .A0(n5323), .A1(n6040), .B0(n4538), .B1(n5668), .C0(n5242), 
        .C1(n5990), .Y(n5667) );
  AOI221XL U6688 ( .A0(n5331), .A1(n5997), .B0(n5333), .B1(n6039), .C0(n5669), 
        .Y(n5668) );
  OAI22XL U6689 ( .A0(n5972), .A1(n4561), .B0(pattern_after[23]), .B1(n4587), 
        .Y(n5669) );
  AOI2BB1X1 U6690 ( .A0N(n4563), .A1N(n5297), .B0(pattern[32]), .Y(n5249) );
  AOI2BB1X1 U6691 ( .A0N(n4568), .A1N(n5309), .B0(pattern[28]), .Y(n5238) );
  AOI2BB1X1 U6692 ( .A0N(n4598), .A1N(n5309), .B0(pattern[30]), .Y(n5239) );
  AOI2BB1X1 U6693 ( .A0N(n4588), .A1N(n5309), .B0(pattern[31]), .Y(n5233) );
  AOI2BB1X1 U6694 ( .A0N(n4599), .A1N(n5297), .B0(pattern[38]), .Y(n5217) );
  AOI2BB1X1 U6695 ( .A0N(n4589), .A1N(n5297), .B0(pattern[39]), .Y(n5218) );
  AOI2BB1X1 U6696 ( .A0N(n4569), .A1N(n5297), .B0(pattern[36]), .Y(n5219) );
  AND2X2 U6697 ( .A(n5427), .B(n5428), .Y(n5405) );
  NOR4X1 U6698 ( .A(pattern[8]), .B(pattern[15]), .C(pattern[14]), .D(
        pattern[12]), .Y(n5428) );
  NOR4X1 U6699 ( .A(n5978), .B(n5984), .C(n5980), .D(n6011), .Y(n5427) );
  AND4X1 U6700 ( .A(pattern[18]), .B(n4555), .C(pattern[21]), .D(n5490), .Y(
        n5385) );
  NOR3X1 U6701 ( .A(pattern[20]), .B(pattern[23]), .C(pattern[22]), .Y(n5490)
         );
  AND4X1 U6702 ( .A(pattern[3]), .B(pattern[2]), .C(n5426), .D(pattern[1]), 
        .Y(n5425) );
  NOR2X1 U6703 ( .A(pattern[7]), .B(pattern[0]), .Y(n5426) );
  NAND4X1 U6704 ( .A(n5768), .B(n5769), .C(n5770), .D(n5771), .Y(n5737) );
  NAND3X1 U6705 ( .A(pattern[17]), .B(n5385), .C(pattern[19]), .Y(n5376) );
  OAI221X1 U6706 ( .A0(n5588), .A1(n5502), .B0(n5589), .B1(n5927), .C0(n5928), 
        .Y(n5111) );
  AOI2BB2X1 U6707 ( .B0(n5521), .B1(n6456), .A0N(n5929), .A1N(n5498), .Y(n5928) );
  OAI22XL U6708 ( .A0(stringData[183]), .A1(n6476), .B0(stringData[247]), .B1(
        n6349), .Y(n5930) );
  AOI222XL U6709 ( .A0(stringData[117]), .A1(n6376), .B0(stringData[181]), 
        .B1(n6359), .C0(stringData[245]), .C1(n6356), .Y(n5509) );
  AOI2BB2X1 U6710 ( .B0(n4863), .B1(n5512), .A0N(n5502), .A1N(n5513), .Y(n5511) );
  AOI222XL U6711 ( .A0(stringData[112]), .A1(n6376), .B0(stringData[176]), 
        .B1(n6359), .C0(stringData[240]), .C1(n6356), .Y(n5497) );
  AOI2BB2X1 U6712 ( .B0(n4863), .B1(n5501), .A0N(n5502), .A1N(n5503), .Y(n5500) );
  AOI222XL U6713 ( .A0(stringData[116]), .A1(n6375), .B0(stringData[180]), 
        .B1(n6359), .C0(stringData[244]), .C1(n6356), .Y(n5504) );
  AOI2BB2X1 U6714 ( .B0(n4863), .B1(n5507), .A0N(n5502), .A1N(n5508), .Y(n5506) );
  NAND4X2 U6715 ( .A(pattern_after[5]), .B(n5730), .C(n6013), .D(n5985), .Y(
        n5695) );
  AOI222XL U6716 ( .A0(stringData[115]), .A1(n6376), .B0(stringData[179]), 
        .B1(n6359), .C0(stringData[243]), .C1(n6356), .Y(n5914) );
  AOI2BB2X1 U6717 ( .B0(n4863), .B1(n5888), .A0N(n5872), .A1N(n5502), .Y(n5915) );
  AOI222XL U6718 ( .A0(stringData[113]), .A1(n6376), .B0(stringData[177]), 
        .B1(n6359), .C0(stringData[241]), .C1(n6356), .Y(n5905) );
  AOI2BB2X1 U6719 ( .B0(n4863), .B1(n5601), .A0N(n5502), .A1N(n5602), .Y(n5906) );
  AOI22X1 U6720 ( .A0(stringData[96]), .A1(n6303), .B0(n5585), .B1(n6468), .Y(
        n5584) );
  AOI22X1 U6721 ( .A0(stringData[99]), .A1(n6303), .B0(n5814), .B1(n6474), .Y(
        n5917) );
  AOI22X1 U6722 ( .A0(stringData[97]), .A1(n6303), .B0(n5775), .B1(n6468), .Y(
        n5908) );
  AOI22X1 U6723 ( .A0(stringData[102]), .A1(n6303), .B0(n5651), .B1(n6468), 
        .Y(n5952) );
  AOI22X1 U6724 ( .A0(stringData[98]), .A1(n6303), .B0(n5828), .B1(n6468), .Y(
        n5942) );
  AOI22X1 U6725 ( .A0(stringData[103]), .A1(n6303), .B0(n5648), .B1(n6474), 
        .Y(n5936) );
  OAI222XL U6726 ( .A0(n5568), .A1(n5999), .B0(n4477), .B1(n5569), .C0(n5570), 
        .C1(n6061), .Y(n5567) );
  AOI221XL U6727 ( .A0(n5257), .A1(n6002), .B0(n5571), .B1(n6054), .C0(n5572), 
        .Y(n5569) );
  OAI22XL U6728 ( .A0(pattern_after[44]), .A1(n4570), .B0(n5973), .B1(n4564), 
        .Y(n5572) );
  OAI222XL U6729 ( .A0(n5608), .A1(n6003), .B0(n4490), .B1(n5609), .C0(n5610), 
        .C1(n6055), .Y(n5607) );
  AOI221XL U6730 ( .A0(n5611), .A1(n6044), .B0(n5612), .B1(n5995), .C0(n5613), 
        .Y(n5609) );
  OAI22XL U6731 ( .A0(pattern_after[38]), .A1(n4599), .B0(pattern_after[39]), 
        .B1(n4589), .Y(n5613) );
  NAND2X1 U6732 ( .A(special), .B(n4516), .Y(n5475) );
  NAND3X2 U6733 ( .A(pattern[25]), .B(n5339), .C(pattern[27]), .Y(n5309) );
  XOR2X1 U6734 ( .A(\sub_1_root_add_0_root_add_92_2/n1 ), .B(n5477), .Y(n5487)
         );
  AOI22X1 U6735 ( .A0(N176), .A1(n5484), .B0(n4515), .B1(N170), .Y(n5488) );
  XOR2X1 U6736 ( .A(\sub_1_root_sub_52_S2_2/carry[3] ), .B(stringNum[3]), .Y(
        n5485) );
  AOI22X1 U6737 ( .A0(N175), .A1(n5484), .B0(N169), .B1(n4515), .Y(n5486) );
  AOI2BB1X1 U6738 ( .A0N(n5167), .A1N(n5111), .B0(pattern[63]), .Y(n5110) );
  AOI2BB1X1 U6739 ( .A0N(n4600), .A1N(n5286), .B0(pattern[46]), .Y(n5205) );
  AOI2BB1X1 U6740 ( .A0N(n4565), .A1N(n5274), .B0(pattern[48]), .Y(n5185) );
  AOI2BB1X1 U6741 ( .A0N(n4596), .A1N(n5274), .B0(pattern[54]), .Y(n5258) );
  AOI2BB1X1 U6742 ( .A0N(n4595), .A1N(n5167), .B0(pattern[62]), .Y(n5108) );
  AOI2BB1X1 U6743 ( .A0N(n4570), .A1N(n5286), .B0(pattern[44]), .Y(n5208) );
  AOI2BB1X1 U6744 ( .A0N(n4564), .A1N(n5286), .B0(pattern[40]), .Y(n5250) );
  AOI2BB1X1 U6745 ( .A0N(n4590), .A1N(n5286), .B0(pattern[47]), .Y(n5200) );
  AOI2BB1X1 U6746 ( .A0N(n4586), .A1N(n5274), .B0(pattern[55]), .Y(n5191) );
  AOI2BB1X1 U6747 ( .A0N(n4571), .A1N(n5274), .B0(pattern[52]), .Y(n5188) );
  AOI2BB1X1 U6748 ( .A0N(n4566), .A1N(n5167), .B0(pattern[56]), .Y(n5118) );
  AOI2BB1X1 U6749 ( .A0N(n4572), .A1N(n5167), .B0(pattern[60]), .Y(n5116) );
  AND4X1 U6750 ( .A(pattern[26]), .B(n4871), .C(pattern[29]), .D(n5492), .Y(
        n5339) );
  NOR3X1 U6751 ( .A(pattern[28]), .B(pattern[31]), .C(pattern[30]), .Y(n5492)
         );
  AND4X1 U6752 ( .A(pattern[34]), .B(n6018), .C(pattern[37]), .D(n5491), .Y(
        n5340) );
  NOR3X1 U6753 ( .A(pattern[36]), .B(pattern[39]), .C(pattern[38]), .Y(n5491)
         );
  AND4X1 U6754 ( .A(pattern[42]), .B(n6019), .C(pattern[45]), .D(n5495), .Y(
        n5341) );
  NOR3X1 U6755 ( .A(pattern[44]), .B(pattern[47]), .C(pattern[46]), .Y(n5495)
         );
  AND4X1 U6756 ( .A(pattern[50]), .B(n6020), .C(pattern[53]), .D(n5494), .Y(
        n5343) );
  NOR3X1 U6757 ( .A(pattern[52]), .B(pattern[55]), .C(pattern[54]), .Y(n5494)
         );
  AND4X1 U6758 ( .A(pattern[58]), .B(n6017), .C(pattern[61]), .D(n5493), .Y(
        n5263) );
  NOR3X1 U6759 ( .A(pattern[60]), .B(pattern[63]), .C(pattern[62]), .Y(n5493)
         );
  NAND4X1 U6760 ( .A(pattern_after[6]), .B(pattern_after[4]), .C(n5730), .D(
        n6014), .Y(n5724) );
  CLKINVX1 U6761 ( .A(n5948), .Y(n4595) );
  OAI221XL U6762 ( .A0(n5949), .A1(n5498), .B0(n6296), .B1(n5532), .C0(n5950), 
        .Y(n5948) );
  AOI222XL U6763 ( .A0(stringData[118]), .A1(n6376), .B0(stringData[182]), 
        .B1(n6359), .C0(stringData[246]), .C1(n6356), .Y(n5949) );
  AOI2BB2X1 U6764 ( .B0(n4863), .B1(n5592), .A0N(n5502), .A1N(n5593), .Y(n5950) );
  CLKINVX1 U6765 ( .A(n5938), .Y(n4591) );
  OAI221XL U6766 ( .A0(n5939), .A1(n5498), .B0(n6296), .B1(n5549), .C0(n5940), 
        .Y(n5938) );
  AOI222XL U6767 ( .A0(stringData[114]), .A1(n6376), .B0(stringData[178]), 
        .B1(n6359), .C0(stringData[242]), .C1(n6356), .Y(n5939) );
  AOI2BB2X1 U6768 ( .B0(n4863), .B1(n5894), .A0N(n5502), .A1N(n5866), .Y(n5940) );
  AND4X1 U6769 ( .A(pattern_after[3]), .B(pattern_after[2]), .C(n5731), .D(
        pattern_after[1]), .Y(n5730) );
  NOR2X1 U6770 ( .A(pattern_after[7]), .B(pattern_after[0]), .Y(n5731) );
  NAND3X1 U6771 ( .A(patternCounter[3]), .B(n6004), .C(n5109), .Y(n5105) );
  XNOR2X1 U6772 ( .A(n5110), .B(n5111), .Y(n5109) );
  XOR2X1 U6773 ( .A(\r685/carry[4] ), .B(\sub_1_root_add_0_root_add_92_2/n1 ), 
        .Y(N170) );
  OAI21X1 U6774 ( .A0(\sub_1_root_add_0_root_add_92_2/n3 ), .A1(n6348), .B0(
        \sub_1_root_add_0_root_add_92_2/carry[1] ), .Y(N166) );
  XNOR2X1 U6775 ( .A(n5481), .B(n6296), .Y(n5387) );
  OAI21XL U6776 ( .A0(n5475), .A1(n5482), .B0(n5483), .Y(n5481) );
  XOR2X1 U6777 ( .A(\sub_1_root_add_0_root_add_92_2/n3 ), .B(n6350), .Y(n5482)
         );
  OAI22XL U6778 ( .A0(N166), .A1(n5484), .B0(n4515), .B1(n4833), .Y(n5483) );
  OAI31XL U6779 ( .A0(n4571), .A1(pattern_after[52]), .A2(n4473), .B0(n5519), 
        .Y(n5516) );
  AOI32X1 U6780 ( .A0(n5261), .A1(n6066), .A2(n5520), .B0(pattern_after[55]), 
        .B1(n4586), .Y(n5519) );
  NAND3X2 U6781 ( .A(pattern[33]), .B(n5340), .C(pattern[35]), .Y(n5297) );
  NAND3X2 U6782 ( .A(pattern[41]), .B(n5341), .C(pattern[43]), .Y(n5286) );
  XOR2X1 U6783 ( .A(stringNum[5]), .B(\add_0_root_add_51/carry[5] ), .Y(n5479)
         );
  XOR2X1 U6784 ( .A(n5476), .B(stringNum[5]), .Y(n5474) );
  XOR2X1 U6785 ( .A(n5478), .B(stringNum[5]), .Y(n5471) );
  XOR2X1 U6786 ( .A(n5478), .B(n5479), .Y(n5473) );
  NAND2X1 U6787 ( .A(\sub_1_root_add_0_root_add_92_2/n3 ), .B(n6348), .Y(
        \sub_1_root_add_0_root_add_92_2/carry[1] ) );
  AND4X1 U6788 ( .A(pattern_after[18]), .B(n5990), .C(pattern_after[21]), .D(
        n5826), .Y(n5825) );
  NOR3X1 U6789 ( .A(pattern_after[20]), .B(pattern_after[23]), .C(
        pattern_after[22]), .Y(n5826) );
  NOR2X1 U6790 ( .A(\sub_1_root_sub_52_S2_2/carry[3] ), .B(stringNum[3]), .Y(
        n5477) );
  NAND2BX1 U6791 ( .AN(\r685/carry[4] ), .B(
        \sub_1_root_add_0_root_add_92_2/n1 ), .Y(n5478) );
  CLKBUFX3 U6792 ( .A(patternCounter[0]), .Y(n6348) );
  NAND2X1 U6793 ( .A(n5477), .B(\sub_1_root_add_0_root_add_92_2/n1 ), .Y(n5476) );
  CLKBUFX3 U6794 ( .A(n589), .Y(n6350) );
  NOR2X1 U6795 ( .A(\sub_1_root_add_0_root_add_92_2/n3 ), .B(n5991), .Y(
        \sub_1_root_sub_52_S2_2/carry[1] ) );
  NAND3X2 U6796 ( .A(pattern[49]), .B(n5343), .C(pattern[51]), .Y(n5274) );
  NAND3X2 U6797 ( .A(pattern[57]), .B(n5263), .C(pattern[59]), .Y(n5167) );
  AND4X1 U6798 ( .A(pattern_after[34]), .B(n5995), .C(pattern_after[37]), .D(
        n5877), .Y(n5876) );
  NOR3X1 U6799 ( .A(pattern_after[36]), .B(pattern_after[39]), .C(
        pattern_after[38]), .Y(n5877) );
  AND4X1 U6800 ( .A(pattern_after[26]), .B(n5993), .C(pattern_after[29]), .D(
        n5856), .Y(n5855) );
  NOR3X1 U6801 ( .A(pattern_after[28]), .B(pattern_after[31]), .C(
        pattern_after[30]), .Y(n5856) );
  NAND4X1 U6802 ( .A(n5968), .B(n5969), .C(n5970), .D(n5971), .Y(n5741) );
  AND4X1 U6803 ( .A(pattern_after[42]), .B(n5999), .C(pattern_after[45]), .D(
        n5904), .Y(n5891) );
  NOR3X1 U6804 ( .A(pattern_after[44]), .B(pattern_after[47]), .C(
        pattern_after[46]), .Y(n5904) );
  NAND3X2 U6805 ( .A(pattern_after[49]), .B(n5553), .C(pattern_after[51]), .Y(
        n5520) );
  XNOR2X1 U6806 ( .A(n5925), .B(patternCounter[3]), .Y(n5435) );
  OAI21XL U6807 ( .A0(n5924), .A1(n5089), .B0(n5090), .Y(n5925) );
  XOR2X1 U6808 ( .A(\sub_1_root_add_0_root_add_92_2/n1 ), .B(
        \sub_1_root_add_0_root_add_92_2/carry[4] ), .Y(n5061) );
  NAND2X1 U6809 ( .A(patternCounter[2]), .B(n6021), .Y(n4976) );
  NOR2X1 U6810 ( .A(n4858), .B(patternCounter[2]), .Y(n5089) );
  NAND2X1 U6811 ( .A(patternCounter[1]), .B(n4859), .Y(n5093) );
  NOR2X1 U6812 ( .A(n4859), .B(patternCounter[1]), .Y(n5092) );
  AND4X1 U6813 ( .A(pattern_after[50]), .B(n6052), .C(pattern_after[53]), .D(
        n5557), .Y(n5553) );
  NOR3X1 U6814 ( .A(pattern_after[52]), .B(pattern_after[55]), .C(
        pattern_after[54]), .Y(n5557) );
  XOR2X1 U6815 ( .A(n5060), .B(stringNum[5]), .Y(n5059) );
  NAND2X1 U6816 ( .A(\add_0_root_add_0_root_add_92_2/carry[4] ), .B(n5061), 
        .Y(n5060) );
  XOR2X1 U6817 ( .A(special_locate[2]), .B(special_locate[1]), .Y(N240) );
  NOR2X1 U6818 ( .A(n6350), .B(n4833), .Y(\add_0_root_add_0_root_add_92_2/n1 )
         );
  NAND2X1 U6819 ( .A(n6348), .B(patternCounter[1]), .Y(n4974) );
  XOR2X1 U6820 ( .A(\sub_1_root_add_0_root_add_92_2/n3 ), .B(n6295), .Y(n5057)
         );
  NAND2X1 U6821 ( .A(special_locate[1]), .B(n6350), .Y(n5079) );
  NAND2X1 U6822 ( .A(special_locate[1]), .B(n5991), .Y(n5076) );
  OR2X1 U6823 ( .A(n6293), .B(\sub_1_root_add_0_root_add_92_2/carry[4] ), .Y(
        n5058) );
  INVX3 U6824 ( .A(n375), .Y(n4849) );
  INVX3 U6825 ( .A(n5977), .Y(n4468) );
  XOR2X1 U6826 ( .A(n5087), .B(patternCounter[3]), .Y(n5038) );
  OAI21XL U6827 ( .A0(n5088), .A1(n5089), .B0(n5090), .Y(n5087) );
  NOR2X1 U6828 ( .A(n6350), .B(n6454), .Y(\add_653_S2/carry[1] ) );
  CLKINVX1 U6829 ( .A(reset), .Y(n4836) );
endmodule

